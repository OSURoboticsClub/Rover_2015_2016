// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Thu Apr  7 00:09:07 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    output expansion4 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire n30467 /* synthesis nomerge= */ ;
    
    wire GND_net, VCC_net, n9970_c, n9969, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, signal_light_c, rc_ch1_c, rc_ch2_c, rc_ch3_c, rc_ch4_c, 
        rc_ch7_c, rc_ch8_c, motor_pwm_l_c, xbee_pause_c, debug_c_7, 
        debug_c_5, debug_c_4, debug_c_3, debug_c_2;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire rw, n13252, n13363;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    
    wire clk_255kHz, n27539, n28430, n32, n24716, n962, n1, n2, 
        n26899, n19, n32_adj_477, n2_adj_478, n1_adj_479, n2_adj_480, 
        n13009;
    wire [7:0]n7684;
    
    wire n22, n1_adj_481, n12995, n12;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n24231, n24230, n24229, n24228, n12981, n24227, n24226, 
        n24225, n1_adj_482, n2736, n17481, n17488, n26439, n26939, 
        n2650, n3539, n26922, n2622, n4, n1_adj_483, n2_adj_484, 
        n8472;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire clk_1Hz, prev_clk_1Hz;
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[12:21])
    
    wire prev_select, n2615;
    wire [7:0]n5062;
    
    wire n24822;
    wire [7:0]\register[1]_adj_725 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]\register[0]_adj_726 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]read_value_adj_727;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(92[12:22])
    wire [2:0]read_size_adj_728;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(93[12:21])
    
    wire n64, n7591;
    wire [15:0]n281;
    
    wire n7, n241, n2610;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched, prev_limit_latched;
    wire [31:0]read_value_adj_735;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_736;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_527, n62, n151;
    wire [3:0]n30602;
    
    wire n12795, n26540;
    wire [31:0]n99_adj_1080;
    
    wire n1_adj_529, n7174, n24744, n26896, n3626, n233, n12781;
    wire [7:0]control_reg_adj_745;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched_adj_531, prev_limit_latched_adj_532, step_clk, 
        prev_step_clk;
    wire [31:0]read_value_adj_748;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_749;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_567, n52, n8336;
    wire [3:0]n16_adj_1097;
    
    wire n8430, n7486, n27505, n27503;
    wire [7:0]n571_adj_766;
    
    wire n27502, n28400, n28399;
    wire [31:0]n580_adj_767;
    
    wire n30468;
    wire [7:0]control_reg_adj_785;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_786;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_787;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched_adj_570, prev_limit_latched_adj_571, int_step, 
        step_clk_adj_572, prev_step_clk_adj_573;
    wire [31:0]read_value_adj_788;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_789;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_608, n7140, n7452, n3356, n3452, n27784, 
        n27783, n27782, n22_adj_609, n32_adj_610, n26512;
    wire [7:0]control_reg_adj_825;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched_adj_612, prev_limit_latched_adj_613;
    wire [31:0]read_value_adj_828;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_829;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_648, n7382, n19316;
    wire [31:0]n580_adj_847;
    
    wire n15, n15_adj_649, n11054, n176, n28582, n18265, n13, 
        n18268, n14, n8273, n28403, n7348, n12650, n12649, n12647, 
        n6, n12605, n12599, n12585, n12583, n12580, n2_adj_650, 
        n26558, n11, n28425, n28576, n2_adj_651, n4_adj_652;
    wire [14:0]n66_adj_1219;
    
    wire n24721, n6_adj_654, n4_adj_655, n1_adj_656, n4_adj_657, n4_adj_658, 
        n27027, n19804, n1_adj_659, n2_adj_660, n1_adj_661, n2_adj_662, 
        n1_adj_663, n2_adj_664, n1_adj_665, n2_adj_666, n1_adj_667, 
        n4_adj_668, n4_adj_669, n4_adj_670, n27025, n2_adj_671, n1_adj_672, 
        n2_adj_673, n1_adj_674, n2_adj_675, n1_adj_676, n2_adj_677, 
        n1_adj_678, n2_adj_679, n1_adj_680, n2_adj_681, n1_adj_682, 
        n2_adj_683, n26514, n26090, n1_adj_684, n2_adj_685, n1_adj_686, 
        n2_adj_687, n1_adj_688, n2_adj_689, n2_adj_690, n1_adj_691, 
        n2_adj_692, n1_adj_693, n2_adj_694, n19338, n28563, n28560, 
        n18270, n18276, n18278, n12_adj_695, n28415, n26556, n26489, 
        n10109, n26396, n13536, n13535, n13534, n28414, n10107, 
        n16717;
    wire [3:0]n6596;
    
    wire n7278, n13527, n26437, n26425, n14714, n14876, n14875, 
        n14873, n28542, n28537, n24707;
    wire [7:0]n7702;
    
    wire n26102, n28402, n26076, n1_adj_696;
    wire [31:0]n6021;
    
    wire n26949, n26947;
    wire [7:0]n7693;
    
    wire n30, n13489, n82;
    wire [3:0]state_adj_885;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    
    wire select_clk, n27040;
    wire [31:0]n59;
    
    wire n28508, n24755, n28506, n26907, n46, n28411, n28505, 
        n28504, n27035, n24633, n28401, n28410, n30_adj_697, n10, 
        n9, n8, n41, n31, n27023, n32_adj_698, n28, n29, n21, 
        n22_adj_699, n28487, n28485, n28482, n28480, n24832, n28477, 
        n28476, n19370, n2_adj_700, n10035, n26087, n4_adj_701, 
        n27504, n26101, n26097, n26089, n26091, n26077, n26078, 
        n26082, n26084, n26099, n26086, n26080, n26088, n7244, 
        n26085, n79_adj_702, n26096, n26094, n26092, n26093, n26081, 
        n7001, n26095, n14_adj_703, n25733, n26079, n26083, n24815, 
        n26103, n26098, n14798, n26100, n24743, n30473, n24741, 
        n6966, n1_adj_704, n24551, n28458, n28457, n30471, n28406, 
        n28405, n28452, n28451, n19865, n30470, n28448, n28445, 
        n28443, n28442, n28441, n28440, n28439, n30469;
    wire [3:0]state_adj_1029;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n28438, n27404, n47, n11943, n26942, n26945, n28431;
    
    VHI i2 (.Z(VCC_net));
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .debug_c_c(debug_c_c), 
            .n12981(n12981), .n28477(n28477), .databus({databus}), .VCC_net(VCC_net), 
            .GND_net(GND_net), .Stepper_Z_nFault_c(Stepper_Z_nFault_c), 
            .\read_size[0] (read_size_adj_789[0]), .n13252(n13252), .n233(n233), 
            .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n12995(n12995), .n579(n571_adj_766[0]), 
            .prev_step_clk(prev_step_clk_adj_573), .step_clk(step_clk_adj_572), 
            .limit_latched(limit_latched_adj_570), .prev_limit_latched(prev_limit_latched_adj_571), 
            .prev_select(prev_select_adj_608), .n28487(n28487), .\read_size[2] (read_size_adj_789[2]), 
            .n26489(n26489), .n28438(n28438), .\div_factor_reg[9] (div_factor_reg_adj_786[9]), 
            .\div_factor_reg[6] (div_factor_reg_adj_786[6]), .\div_factor_reg[5] (div_factor_reg_adj_786[5]), 
            .n608(n580_adj_847[4]), .n610(n580_adj_847[2]), .\control_reg[7] (control_reg_adj_785[7]), 
            .n28445(n28445), .n10109(n10109), .Stepper_Z_En_c(Stepper_Z_En_c), 
            .Stepper_Z_Dir_c(Stepper_Z_Dir_c), .\control_reg[3] (control_reg_adj_785[3]), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), 
            .read_value({read_value_adj_788}), .n3452(n3452), .\steps_reg[9] (steps_reg_adj_787[9]), 
            .\steps_reg[5] (steps_reg_adj_787[5]), .\steps_reg[6] (steps_reg_adj_787[6]), 
            .\steps_reg[3] (steps_reg_adj_787[3]), .n32(n32_adj_477), .limit_c_2(limit_c_2), 
            .n24832(n24832), .n6050(n6021[3]), .n18278(n18278), .n18270(n18270), 
            .n79(n99_adj_1080[9]), .int_step(int_step), .n22(n22), .n28410(n28410), 
            .\div_factor_reg[3] (div_factor_reg_adj_786[3]), .n7694(n7693[7]), 
            .n28402(n28402), .n14875(n14875), .n7382(n7382), .n7348(n7348)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(588[25] 601[45])
    LUT4 i8_2_lut (.A(state_adj_885[1]), .B(state_adj_885[0]), .Z(n6596[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    defparam i8_2_lut.init = 16'h6666;
    LUT4 i1_4_lut (.A(n28477), .B(n46), .C(state_adj_1029[3]), .D(state_adj_1029[2]), 
         .Z(n30602[2])) /* synthesis lut_function=(!(A+(B (D)+!B (C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0144;
    LUT4 i1_2_lut_rep_284_3_lut_3_lut_4_lut (.A(n82), .B(reset_count[14]), 
         .C(n7591), .D(select_clk), .Z(n28405)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_284_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i13337_2_lut_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(databus[0]), 
         .Z(n571_adj_766[0])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13337_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(n28487), .D(prev_select_adj_608), 
         .Z(n13252)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(n8273), .Z(n13363)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_adj_401 (.A(n82), .B(reset_count[14]), .C(n12649), 
         .Z(n12650)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_401.init = 16'hf7f7;
    LUT4 i1_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(n151), .D(n28482), 
         .Z(n2622)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0800;
    LUT4 state_1__bdd_4_lut_20573 (.A(state_adj_1029[1]), .B(state_adj_1029[3]), 
         .C(state_adj_1029[2]), .D(state_adj_1029[0]), .Z(n27404)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)+!B !(C+(D))))) */ ;
    defparam state_1__bdd_4_lut_20573.init = 16'h373e;
    LUT4 i925_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(select[1]), 
         .D(prev_select), .Z(n12585)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i925_3_lut_4_lut.init = 16'h0080;
    LUT4 i2450_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(clk_1Hz), 
         .D(prev_clk_1Hz), .Z(n8430)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i2450_3_lut_4_lut.init = 16'h77f7;
    LUT4 i13532_2_lut_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(databus[1]), 
         .Z(n580_adj_767[1])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13532_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i4036_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(limit_latched), 
         .D(prev_limit_latched), .Z(n10035)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i4036_3_lut_4_lut.init = 16'h77f7;
    LUT4 i8870_2_lut_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(n7382), 
         .D(n7348), .Z(n14875)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i8870_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1_2_lut_3_lut_adj_402 (.A(n82), .B(reset_count[14]), .C(n12580), 
         .Z(n12583)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_402.init = 16'hf7f7;
    LUT4 i2_3_lut_4_lut_adj_403 (.A(n82), .B(reset_count[14]), .C(n28480), 
         .D(prev_select_adj_527), .Z(n2615)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut_adj_403.init = 16'h0080;
    LUT4 i13482_2_lut_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(databus[7]), 
         .Z(n281[15])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13482_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i988_2_lut_rep_281_3_lut (.A(n82), .B(reset_count[14]), .C(n7348), 
         .Z(n28402)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i988_2_lut_rep_281_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_309_3_lut (.A(n82), .B(reset_count[14]), .C(prev_select_adj_648), 
         .Z(n28430)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_309_3_lut.init = 16'h0808;
    LUT4 i2_3_lut_rep_464 (.A(n82), .B(reset_count[14]), .C(n6966), .D(clk_255kHz), 
         .Z(n30469)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_464.init = 16'h0080;
    LUT4 i2_3_lut_rep_465 (.A(n82), .B(reset_count[14]), .C(n6966), .D(clk_255kHz), 
         .Z(n30470)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_465.init = 16'h0080;
    LUT4 i13392_2_lut (.A(reset_count[9]), .B(reset_count[10]), .Z(n19370)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13392_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_rep_466 (.A(n82), .B(reset_count[14]), .C(n6966), .D(clk_255kHz), 
         .Z(n30471)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_466.init = 16'h0080;
    LUT4 i13928_4_lut_rep_364 (.A(reset_count[12]), .B(reset_count[14]), 
         .C(reset_count[13]), .D(n26512), .Z(n28485)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i13928_4_lut_rep_364.init = 16'hfcec;
    LUT4 i13953_1_lut_rep_336_4_lut (.A(reset_count[12]), .B(reset_count[14]), 
         .C(reset_count[13]), .D(n26512), .Z(n28457)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C (D))))) */ ;
    defparam i13953_1_lut_rep_336_4_lut.init = 16'h0313;
    LUT4 i13953_1_lut_rep_468 (.A(reset_count[12]), .B(reset_count[14]), 
         .C(reset_count[13]), .D(n26512), .Z(n30473)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C (D))))) */ ;
    defparam i13953_1_lut_rep_468.init = 16'h0313;
    LUT4 state_1__bdd_4_lut (.A(state_adj_1029[1]), .B(state_adj_1029[0]), 
         .C(n962), .D(state_adj_1029[3]), .Z(n27539)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h7ffe;
    PFUMX i10746 (.BLUT(n59[2]), .ALUT(n32_adj_698), .C0(n7), .Z(n5062[2]));
    PFUMX i10741 (.BLUT(n59[4]), .ALUT(n31), .C0(n7), .Z(n5062[4]));
    PFUMX i10736 (.BLUT(n59[5]), .ALUT(n30_adj_697), .C0(n7), .Z(n5062[5]));
    PFUMX i10731 (.BLUT(n59[3]), .ALUT(n29), .C0(n7), .Z(n5062[3]));
    PFUMX i10726 (.BLUT(n22_adj_699), .ALUT(n28), .C0(n7), .Z(n5062[1]));
    FD1P3AX reset_count_2368_2369__i1 (.D(n66_adj_1219[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i1.GSR = "ENABLED";
    PFUMX i20646 (.BLUT(n27783), .ALUT(n27782), .C0(state_adj_1029[2]), 
          .Z(n27784));
    LUT4 i12292_3_lut (.A(Stepper_Z_Dir_c), .B(div_factor_reg_adj_786[5]), 
         .C(register_addr[1]), .Z(n18276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i12292_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_404 (.A(register_addr[1]), .B(div_factor_reg_adj_786[9]), 
         .C(steps_reg_adj_787[9]), .D(register_addr[0]), .Z(n99_adj_1080[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_404.init = 16'ha088;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    IB n9970_pad (.I(uart_rx), .O(n9970_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    OB debug_pad_0 (.I(n9970_c), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_1 (.I(n9969), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_6 (.I(n28477), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB motor_pwm_r_pad (.I(GND_net), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    OB expansion5_pad (.I(GND_net), .O(expansion5));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    OB expansion4_pad (.I(GND_net), .O(expansion4));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    OB expansion3_pad (.I(GND_net), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    OB expansion2_pad (.I(GND_net), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion1_pad (.I(GND_net), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    LUT4 i12284_3_lut (.A(Stepper_Z_En_c), .B(div_factor_reg_adj_786[6]), 
         .C(register_addr[1]), .Z(n18268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i12284_3_lut.init = 16'hcaca;
    LUT4 i12281_3_lut (.A(control_reg_adj_785[3]), .B(div_factor_reg_adj_786[3]), 
         .C(register_addr[1]), .Z(n18265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i12281_3_lut.init = 16'hcaca;
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB uart_tx_pad (.I(n9969), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    LUT4 i1_4_lut_adj_405 (.A(n41), .B(n28508), .C(n17488), .D(n28443), 
         .Z(n21)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_405.init = 16'h5154;
    LUT4 state_3__bdd_4_lut (.A(state_adj_1029[3]), .B(state_adj_1029[1]), 
         .C(state_adj_1029[0]), .D(n962), .Z(n27783)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam state_3__bdd_4_lut.init = 16'h8f0e;
    LUT4 state_3__bdd_2_lut (.A(state_adj_1029[3]), .B(state_adj_1029[0]), 
         .Z(n27782)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_3__bdd_2_lut.init = 16'h1111;
    LUT4 m1_lut (.Z(n30467)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    LUT4 i1_4_lut_adj_406 (.A(n41), .B(\register[0]_adj_726 [1]), .C(n14_adj_703), 
         .D(n28537), .Z(n25733)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_406.init = 16'h5051;
    LUT4 i1_4_lut_adj_407 (.A(n17481), .B(n28560), .C(n28537), .D(n4_adj_701), 
         .Z(n14_adj_703)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_407.init = 16'ha8a0;
    LUT4 i20432_4_lut (.A(reset_count[14]), .B(n79_adj_702), .C(n19370), 
         .D(n26558), .Z(n30)) /* synthesis lut_function=(!(A (B+(C (D))))) */ ;
    defparam i20432_4_lut.init = 16'h5777;
    LUT4 i1_4_lut_adj_408 (.A(n19804), .B(n26556), .C(reset_count[6]), 
         .D(reset_count[5]), .Z(n26558)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[17:42])
    defparam i1_4_lut_adj_408.init = 16'hfcec;
    LUT4 i13822_4_lut (.A(reset_count[0]), .B(reset_count[4]), .C(n6), 
         .D(reset_count[3]), .Z(n19804)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i13822_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(reset_count[1]), .B(reset_count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(reset_count[11]), .B(reset_count[12]), .C(reset_count[13]), 
         .Z(n79_adj_702)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i2_3_lut.init = 16'hfefe;
    FD1P3AX reset_count_2368_2369__i2 (.D(n66_adj_1219[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i2.GSR = "ENABLED";
    LUT4 i20293_2_lut (.A(int_step), .B(control_reg_adj_785[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i20293_2_lut.init = 16'h9999;
    FD1P3AX reset_count_2368_2369__i3 (.D(n66_adj_1219[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i4 (.D(n66_adj_1219[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i5 (.D(n66_adj_1219[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i6 (.D(n66_adj_1219[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i7 (.D(n66_adj_1219[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i8 (.D(n66_adj_1219[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i9 (.D(n66_adj_1219[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i10 (.D(n66_adj_1219[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i11 (.D(n66_adj_1219[10]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i12 (.D(n66_adj_1219[11]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i13 (.D(n66_adj_1219[12]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i14 (.D(n66_adj_1219[13]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2368_2369__i15 (.D(n66_adj_1219[14]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369__i15.GSR = "ENABLED";
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 i20420_2_lut_rep_356 (.A(n82), .B(reset_count[14]), .Z(n28477)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i20420_2_lut_rep_356.init = 16'h7777;
    LUT4 i980_2_lut_rep_280_3_lut (.A(n82), .B(reset_count[14]), .C(n7140), 
         .Z(n28401)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i980_2_lut_rep_280_3_lut.init = 16'hf7f7;
    LUT4 i2_4_lut (.A(state_adj_1029[3]), .B(n28477), .C(state_adj_1029[2]), 
         .D(n46), .Z(n24633)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam i2_4_lut.init = 16'h1202;
    LUT4 i8743_2_lut_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(n7174), 
         .D(n7140), .Z(n14714)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i8743_2_lut_3_lut_4_lut.init = 16'hf070;
    GlobalControlPeripheral global_control (.debug_c_c(debug_c_c), .n8430(n8430), 
            .n28477(n28477), .read_size({read_size}), .n12585(n12585), 
            .n19316(n19316), .prev_clk_1Hz(prev_clk_1Hz), .clk_1Hz(clk_1Hz), 
            .prev_select(prev_select), .\select[1] (select[1]), .xbee_pause_c(xbee_pause_c), 
            .n28537(n28537), .\register[1][1] (\register[1]_adj_725 [1]), 
            .n28504(n28504), .\control_reg[7] (control_reg_adj_745[7]), 
            .n24822(n24822), .n32(n32_adj_610), .\control_reg[7]_adj_238 (control_reg[7]), 
            .n24815(n24815), .n19(n19), .\register[0][7] (\register[0]_adj_726 [7]), 
            .n28508(n28508), .n19865(n19865), .n28505(n28505), .\register[1][7] (\register[1]_adj_725 [7]), 
            .n28506(n28506), .n19338(n19338), .\register[0][4] (\register[0]_adj_726 [4]), 
            .n17481(n17481), .\control_reg[7]_adj_239 (control_reg_adj_825[7]), 
            .n24744(n24744), .n32_adj_240(n32), .\register[2][31] (\register[2] [31]), 
            .\register[2][30] (\register[2] [30]), .\register[2][29] (\register[2] [29]), 
            .\register[2][28] (\register[2] [28]), .\register[2][27] (\register[2] [27]), 
            .\register[2][26] (\register[2] [26]), .\register[2][25] (\register[2] [25]), 
            .\register[2][24] (\register[2] [24]), .\register[2][23] (\register[2] [23]), 
            .\register[2][22] (\register[2] [22]), .\register[2][21] (\register[2] [21]), 
            .\register[2][20] (\register[2] [20]), .\register[2][19] (\register[2] [19]), 
            .\register[2][18] (\register[2] [18]), .\register[2][17] (\register[2] [17]), 
            .\register[2][16] (\register[2] [16]), .\register[2][15] (\register[2] [15]), 
            .\register[2][14] (\register[2] [14]), .\register[2][13] (\register[2] [13]), 
            .\register[2][12] (\register[2] [12]), .\register[2][11] (\register[2] [11]), 
            .\register[2][10] (\register[2] [10]), .\register[2][9] (\register[2] [9]), 
            .\register[2][8] (\register[2] [8]), .\register[2][7] (\register[2] [7]), 
            .\register[2][6] (\register[2] [6]), .\register[2][5] (\register[2] [5]), 
            .\register[2][4] (\register[2] [4]), .\control_reg[7]_adj_241 (control_reg_adj_785[7]), 
            .n24832(n24832), .n32_adj_242(n32_adj_477), .signal_light_c(signal_light_c), 
            .\register_addr[1] (register_addr[1]), .\register_addr[0] (register_addr[0]), 
            .n27504(n27504), .n27502(n27502), .n11(n11), .n28431(n28431), 
            .rw(rw), .n15(n15_adj_649), .n28582(n28582), .n6(n6_adj_654), 
            .\read_value[2] (read_value[2]), .n27505(n27505), .n27503(n27503), 
            .\read_value[3] (read_value[3]), .n8472(n8472), .\read_value[4] (read_value[4]), 
            .n26100(n26100), .\read_value[5] (read_value[5]), .n26096(n26096), 
            .\read_value[6] (read_value[6]), .n26088(n26088), .\read_value[7] (read_value[7]), 
            .n26090(n26090), .\read_value[8] (read_value[8]), .n26076(n26076), 
            .\read_value[9] (read_value[9]), .n26077(n26077), .\read_value[10] (read_value[10]), 
            .n26081(n26081), .\read_value[11] (read_value[11]), .n26083(n26083), 
            .\read_value[12] (read_value[12]), .n26098(n26098), .\read_value[13] (read_value[13]), 
            .n26085(n26085), .\read_value[14] (read_value[14]), .n26079(n26079), 
            .\read_value[15] (read_value[15]), .n26087(n26087), .\read_value[16] (read_value[16]), 
            .n26084(n26084), .\read_value[17] (read_value[17]), .n26094(n26094), 
            .\read_value[18] (read_value[18]), .n26095(n26095), .\read_value[19] (read_value[19]), 
            .n26093(n26093), .\read_value[20] (read_value[20]), .n26091(n26091), 
            .\read_value[21] (read_value[21]), .n26092(n26092), .\read_value[22] (read_value[22]), 
            .n26080(n26080), .\read_value[23] (read_value[23]), .n26086(n26086), 
            .\read_value[24] (read_value[24]), .n26078(n26078), .\read_value[25] (read_value[25]), 
            .n26082(n26082), .\read_value[26] (read_value[26]), .n26089(n26089), 
            .\read_value[27] (read_value[27]), .n26102(n26102), .\read_value[28] (read_value[28]), 
            .n26097(n26097), .\read_value[29] (read_value[29]), .n26099(n26099), 
            .\read_value[30] (read_value[30]), .n26103(n26103), .\read_value[31] (read_value[31]), 
            .n26101(n26101), .\databus[1] (databus[1]), .GND_net(GND_net), 
            .n26425(n26425), .n62(n62), .n14798(n14798), .n15_adj_243(n15), 
            .\read_value[0] (read_value[0]), .n4(n4), .n2650(n2650), .n26899(n26899)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(495[45] 505[74])
    LUT4 i2_3_lut_rep_282_4_lut (.A(n82), .B(reset_count[14]), .C(n6966), 
         .D(clk_255kHz), .Z(n28403)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_282_4_lut.init = 16'h0080;
    LUT4 i13104_2_lut_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(n6966), 
         .Z(n241)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13104_2_lut_2_lut_3_lut.init = 16'h8080;
    SabertoothSerialPeripheral motor_serial (.\register[1] ({\register[1]_adj_725 [7], 
            Open_0, Open_1, Open_2, Open_3, Open_4, Open_5, Open_6}), 
            .debug_c_c(debug_c_c), .n282(n281[15]), .n28477(n28477), .\databus[6] (databus[6]), 
            .\databus[5] (databus[5]), .\databus[4] (databus[4]), .\databus[3] (databus[3]), 
            .\databus[2] (databus[2]), .\register[1][1] (\register[1]_adj_725 [1]), 
            .\databus[1] (databus[1]), .\databus[0] (databus[0]), .\register[0] ({\register[0]_adj_726 [7], 
            Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, Open_13}), 
            .\register[0][4] (\register[0]_adj_726 [4]), .\register[0][1] (\register[0]_adj_726 [1]), 
            .\read_size[0] (read_size_adj_728[0]), .n28425(n28425), .\select[2] (select[2]), 
            .read_value({read_value_adj_727}), .rw(rw), .n64(n64), .n28415(n28415), 
            .\register_addr[0] (register_addr[0]), .n28560(n28560), .n4(n4_adj_701), 
            .n28537(n28537), .n19865(n19865), .n22(n22_adj_699), .\reset_count[14] (reset_count[14]), 
            .n82(n82), .\register_addr[2] (register_addr[2]), .n28440(n28440), 
            .n28443(n28443), .\state[0] (state_adj_885[0]), .GND_net(GND_net), 
            .n12(n16_adj_1097[0]), .\state[1] (state_adj_885[1]), .n28405(n28405), 
            .n6599(n6596[1]), .n17488(n17488), .n21(n21), .n7(n7), .n19338(n19338), 
            .n25733(n25733), .n28505(n28505), .n962(n962), .n17481(n17481), 
            .n89(n59[2]), .n41(n41), .n32(n32_adj_698), .n87(n59[4]), 
            .n31(n31), .n86(n59[5]), .n30(n30_adj_697), .n88(n59[3]), 
            .n29(n29), .n28(n28), .n5069(n5062[1]), .n5068(n5062[2]), 
            .n5067(n5062[3]), .n5066(n5062[4]), .n5065(n5062[5]), .n28504(n28504), 
            .n28506(n28506), .state({state_adj_1029}), .n27784(n27784), 
            .n13009(n13009), .n24633(n24633), .n19370(n19370), .\reset_count[11] (reset_count[11]), 
            .\reset_count[8] (reset_count[8]), .n24551(n24551), .n26512(n26512), 
            .\reset_count[7] (reset_count[7]), .n26556(n26556), .motor_pwm_l_c(motor_pwm_l_c), 
            .n27404(n27404), .n46(n46), .n7_adj_237(n30602[2]), .\reset_count[6] (reset_count[6]), 
            .\reset_count[5] (reset_count[5]), .\reset_count[4] (reset_count[4]), 
            .n47(n47), .n2736(n2736), .select_clk(select_clk), .n16717(n16717), 
            .n7591(n7591), .n28406(n28406), .n26896(n26896)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(508[29] 516[56])
    LUT4 i1_3_lut_4_lut_4_lut_3_lut_4_lut (.A(n82), .B(reset_count[14]), 
         .C(n28406), .D(state_adj_885[0]), .Z(n16_adj_1097[0])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i1_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2_3_lut_4_lut_adj_409 (.A(n82), .B(reset_count[14]), .C(n27539), 
         .D(state_adj_1029[2]), .Z(n13009)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i2_3_lut_4_lut_adj_409.init = 16'hfff7;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(n26396), 
         .D(n28542), .Z(n12781)) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf777;
    LUT4 i13117_2_lut_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(databus[4]), 
         .Z(n580_adj_847[4])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13117_2_lut_2_lut_3_lut.init = 16'h8080;
    \ProtocolInterface(baud_div=12)  protocol_interface (.register_addr({Open_14, 
            Open_15, Open_16, Open_17, Open_18, register_addr[2:0]}), 
            .n11(n11), .n12585(n12585), .n26425(n26425), .n19316(n19316), 
            .rw(rw), .n28415(n28415), .debug_c_c(debug_c_c), .n30473(n30473), 
            .n28485(n28485), .databus_out({databus_out}), .\select[7] (select[7]), 
            .debug_c_2(debug_c_2), .\select[2] (select[2]), .n28457(n28457), 
            .\select[1] (select[1]), .n28542(n28542), .n28438(n28438), 
            .n26396(n26396), .n28441(n28441), .prev_select(prev_select_adj_567), 
            .n28477(n28477), .n3539(n3539), .\sendcount[1] (sendcount[1]), 
            .n30468(n30468), .databus({databus}), .\read_value[5] (read_value_adj_735[5]), 
            .n4(n4_adj_668), .\read_value[7] (read_value_adj_735[7]), .n4_adj_147(n4_adj_670), 
            .\read_value[0] (read_value_adj_735[0]), .n4_adj_148(n4_adj_652), 
            .\read_value[3] (read_value_adj_735[3]), .n4_adj_149(n4_adj_657), 
            .\read_value[2] (read_value_adj_735[2]), .n4_adj_150(n4_adj_655), 
            .\read_value[4] (read_value_adj_735[4]), .n4_adj_151(n4_adj_658), 
            .n8(n8), .\read_size[0] (read_size_adj_736[0]), .\read_value[6] (read_value_adj_735[6]), 
            .n4_adj_152(n4_adj_669), .n52(n52), .\read_value[13] (read_value_adj_788[13]), 
            .n2(n2_adj_673), .\read_value[10] (read_value_adj_788[10]), 
            .n2_adj_153(n2_adj_660), .\read_value[26] (read_value_adj_788[26]), 
            .n2_adj_154(n2_adj_484), .\read_value[31] (read_value_adj_788[31]), 
            .n2_adj_155(n2_adj_651), .\read_value[29] (read_value_adj_788[29]), 
            .n2_adj_156(n2_adj_700), .\read_value[9] (read_value_adj_788[9]), 
            .n2_adj_157(n2_adj_666), .\read_value[11] (read_value_adj_788[11]), 
            .n2_adj_158(n2_adj_664), .\read_value[30] (read_value_adj_788[30]), 
            .n2_adj_159(n2_adj_650), .\read_value[28] (read_value_adj_788[28]), 
            .n2_adj_160(n2_adj_478), .\read_value[27] (read_value_adj_788[27]), 
            .n2_adj_161(n2_adj_690), .\read_value[25] (read_value_adj_788[25]), 
            .n2_adj_162(n2_adj_480), .\read_value[24] (read_value_adj_788[24]), 
            .n2_adj_163(n2), .\read_value[23] (read_value_adj_788[23]), 
            .n2_adj_164(n2_adj_694), .\read_value[22] (read_value_adj_788[22]), 
            .n2_adj_165(n2_adj_692), .\read_value[21] (read_value_adj_788[21]), 
            .n2_adj_166(n2_adj_685), .\read_value[20] (read_value_adj_788[20]), 
            .n2_adj_167(n2_adj_681), .\read_value[19] (read_value_adj_788[19]), 
            .n2_adj_168(n2_adj_677), .\read_value[18] (read_value_adj_788[18]), 
            .n2_adj_169(n2_adj_683), .\read_value[17] (read_value_adj_788[17]), 
            .n2_adj_170(n2_adj_679), .\read_value[16] (read_value_adj_788[16]), 
            .n2_adj_171(n2_adj_689), .\read_value[15] (read_value_adj_788[15]), 
            .n2_adj_172(n2_adj_687), .\read_value[14] (read_value_adj_788[14]), 
            .n2_adj_173(n2_adj_675), .\read_value[12] (read_value_adj_788[12]), 
            .n2_adj_174(n2_adj_671), .n11943(n11943), .n28563(n28563), 
            .\read_value[8] (read_value_adj_788[8]), .n2_adj_175(n2_adj_662), 
            .n28442(n28442), .n9(n9), .n10(n10), .debug_c_7(debug_c_7), 
            .\reg_size[2] (reg_size[2]), .n28576(n28576), .n28431(n28431), 
            .prev_select_adj_176(prev_select_adj_527), .n28414(n28414), 
            .n28482(n28482), .n151(n151), .n12649(n12649), .n28430(n28430), 
            .n3356(n3356), .prev_select_adj_177(prev_select_adj_608), .n30467(n30467), 
            .\read_value[23]_adj_178 (read_value_adj_828[23]), .n1(n1_adj_693), 
            .\read_value[22]_adj_179 (read_value_adj_828[22]), .n1_adj_180(n1_adj_691), 
            .n26540(n26540), .n8273(n8273), .n3452(n3452), .debug_c_3(debug_c_3), 
            .\register[2][14] (\register[2] [14]), .n26079(n26079), .\register[2][12] (\register[2] [12]), 
            .n26098(n26098), .\register[2][10] (\register[2] [10]), .n26081(n26081), 
            .\register[2][7] (\register[2] [7]), .n26090(n26090), .\register[2][11] (\register[2] [11]), 
            .n26083(n26083), .n28448(n28448), .n28452(n28452), .\control_reg[7] (control_reg_adj_745[7]), 
            .n7685(n7684[7]), .\control_reg[7]_adj_181 (control_reg_adj_785[7]), 
            .n7694(n7693[7]), .\register[2][6] (\register[2] [6]), .n26088(n26088), 
            .\register[2][5] (\register[2] [5]), .n26096(n26096), .\register[2][9] (\register[2] [9]), 
            .n26077(n26077), .\register[2][8] (\register[2] [8]), .n26076(n26076), 
            .\register[2][13] (\register[2] [13]), .n26085(n26085), .\register[2][4] (\register[2] [4]), 
            .n26100(n26100), .n28440(n28440), .n14798(n14798), .n26514(n26514), 
            .\register[2][15] (\register[2] [15]), .n26087(n26087), .\control_reg[7]_adj_182 (control_reg_adj_825[7]), 
            .n7703(n7702[7]), .n28451(n28451), .\register[2][16] (\register[2] [16]), 
            .n26084(n26084), .\register[2][17] (\register[2] [17]), .n26094(n26094), 
            .\register[2][18] (\register[2] [18]), .n26095(n26095), .\steps_reg[5] (steps_reg_adj_787[5]), 
            .n14(n14), .\register[2][19] (\register[2] [19]), .n26093(n26093), 
            .\register[2][20] (\register[2] [20]), .n26091(n26091), .\register[2][21] (\register[2] [21]), 
            .n26092(n26092), .\read_value[21]_adj_183 (read_value_adj_828[21]), 
            .n1_adj_184(n1_adj_684), .n28480(n28480), .\register[2][22] (\register[2] [22]), 
            .n26080(n26080), .\register[2][23] (\register[2] [23]), .n26086(n26086), 
            .n28458(n28458), .\register[2][24] (\register[2] [24]), .n26078(n26078), 
            .\register[2][25] (\register[2] [25]), .n26082(n26082), .\register[2][26] (\register[2] [26]), 
            .n26089(n26089), .\register[2][27] (\register[2] [27]), .n26102(n26102), 
            .\register[2][28] (\register[2] [28]), .n26097(n26097), .\register[2][29] (\register[2] [29]), 
            .n26099(n26099), .\register[2][30] (\register[2] [30]), .n26103(n26103), 
            .n3626(n3626), .n26489(n26489), .n28476(n28476), .n28487(n28487), 
            .n26437(n26437), .n26439(n26439), .n233(n233), .\register[2][31] (\register[2] [31]), 
            .n26101(n26101), .prev_select_adj_185(prev_select_adj_648), 
            .n8472(n8472), .\steps_reg[6] (steps_reg_adj_787[6]), .n13(n13), 
            .\steps_reg[3] (steps_reg_adj_787[3]), .n12(n12_adj_695), .\read_value[20]_adj_186 (read_value_adj_828[20]), 
            .n1_adj_187(n1_adj_680), .debug_c_4(debug_c_4), .\read_value[19]_adj_188 (read_value_adj_828[19]), 
            .n1_adj_189(n1_adj_676), .\read_value[18]_adj_190 (read_value_adj_828[18]), 
            .n1_adj_191(n1_adj_682), .\read_value[17]_adj_192 (read_value_adj_828[17]), 
            .n1_adj_193(n1_adj_678), .n12981(n12981), .\read_value[16]_adj_194 (read_value_adj_828[16]), 
            .n1_adj_195(n1_adj_688), .n15(n15_adj_649), .n8336(n8336), 
            .n4_adj_196(n4), .n12580(n12580), .n62(n62), .n15_adj_197(n15), 
            .n27504(n27504), .n27505(n27505), .n27502(n27502), .n27503(n27503), 
            .n28425(n28425), .n28439(n28439), .n176(n176), .\read_value[15]_adj_198 (read_value_adj_828[15]), 
            .n1_adj_199(n1_adj_686), .debug_c_5(debug_c_5), .\read_value[14]_adj_200 (read_value_adj_828[14]), 
            .n1_adj_201(n1_adj_674), .\read_value[12]_adj_202 (read_value_adj_828[12]), 
            .n1_adj_203(n1_adj_667), .\read_value[8]_adj_204 (read_value_adj_828[8]), 
            .n1_adj_205(n1_adj_661), .n12647(n12647), .\read_value[10]_adj_206 (read_value_adj_828[10]), 
            .n1_adj_207(n1_adj_659), .\read_value[30]_adj_208 (read_value_adj_828[30]), 
            .n1_adj_209(n1_adj_481), .n12599(n12599), .\read_value[9]_adj_210 (read_value_adj_828[9]), 
            .n1_adj_211(n1_adj_665), .\read_value[11]_adj_212 (read_value_adj_828[11]), 
            .n1_adj_213(n1_adj_663), .\read_value[13]_adj_214 (read_value_adj_828[13]), 
            .n1_adj_215(n1_adj_672), .n28445(n28445), .\read_value[27]_adj_216 (read_value_adj_828[27]), 
            .n1_adj_217(n1_adj_696), .\read_value[28]_adj_218 (read_value_adj_828[28]), 
            .n1_adj_219(n1_adj_704), .\read_value[31]_adj_220 (read_value_adj_828[31]), 
            .n1_adj_221(n1_adj_482), .\read_value[29]_adj_222 (read_value_adj_828[29]), 
            .n1_adj_223(n1_adj_529), .\read_value[1] (read_value_adj_828[1]), 
            .n1_adj_224(n1_adj_656), .\read_value[26]_adj_225 (read_value_adj_828[26]), 
            .n1_adj_226(n1_adj_483), .n12995(n12995), .\read_value[25]_adj_227 (read_value_adj_828[25]), 
            .n1_adj_228(n1_adj_479), .\read_value[24]_adj_229 (read_value_adj_828[24]), 
            .n1_adj_230(n1), .\steps_reg[7] (steps_reg[7]), .n12_adj_231(n12), 
            .\reset_count[7] (reset_count[7]), .\reset_count[6] (reset_count[6]), 
            .\reset_count[5] (reset_count[5]), .n24551(n24551), .n9969(n9969), 
            .GND_net(GND_net), .n9970_c(n9970_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[26] 485[57])
    LUT4 i13503_2_lut_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(databus[2]), 
         .Z(n580_adj_847[2])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13503_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i8868_2_lut_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(n7278), 
         .D(n7244), .Z(n14873)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i8868_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i4109_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(limit_latched_adj_570), 
         .D(prev_limit_latched_adj_571), .Z(n10109)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i4109_3_lut_4_lut.init = 16'h77f7;
    LUT4 i984_2_lut_rep_279_3_lut (.A(n82), .B(reset_count[14]), .C(n7244), 
         .Z(n28400)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i984_2_lut_rep_279_3_lut.init = 16'hf7f7;
    LUT4 i992_2_lut_rep_278_3_lut (.A(n82), .B(reset_count[14]), .C(n7452), 
         .Z(n28399)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i992_2_lut_rep_278_3_lut.init = 16'hf7f7;
    LUT4 i8871_2_lut_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(n7486), 
         .D(n7452), .Z(n14876)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i8871_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(n7591), 
         .Z(n16717)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i4107_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(limit_latched_adj_612), 
         .D(prev_limit_latched_adj_613), .Z(n10107)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i4107_3_lut_4_lut.init = 16'h77f7;
    LUT4 i5054_3_lut_4_lut (.A(n82), .B(reset_count[14]), .C(limit_latched_adj_531), 
         .D(prev_limit_latched_adj_532), .Z(n11054)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i5054_3_lut_4_lut.init = 16'h77f7;
    LUT4 i1_2_lut_3_lut_4_lut_adj_410 (.A(n82), .B(reset_count[14]), .C(n26396), 
         .D(n28563), .Z(n12795)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_410.init = 16'h77f7;
    VLO i1 (.Z(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i20299_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(n26896), 
         .Z(n2736)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i20299_2_lut_3_lut.init = 16'hf7f7;
    CCU2D reset_count_2368_2369_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24231), .S0(n66_adj_1219[13]), 
          .S1(n66_adj_1219[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2368_2369_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24230), .COUT(n24231), .S0(n66_adj_1219[11]), 
          .S1(n66_adj_1219[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2368_2369_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24229), .COUT(n24230), .S0(n66_adj_1219[9]), 
          .S1(n66_adj_1219[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2368_2369_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24228), .COUT(n24229), .S0(n66_adj_1219[7]), 
          .S1(n66_adj_1219[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2368_2369_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24227), .COUT(n24228), .S0(n66_adj_1219[5]), 
          .S1(n66_adj_1219[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_7.INJECT1_1 = "NO";
    CCU2D reset_count_2368_2369_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24226), .COUT(n24227), .S0(n66_adj_1219[3]), 
          .S1(n66_adj_1219[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_5.INJECT1_1 = "NO";
    CCU2D reset_count_2368_2369_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24225), .COUT(n24226), .S0(n66_adj_1219[1]), 
          .S1(n66_adj_1219[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2368_2369_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2368_2369_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24225), .S1(n66_adj_1219[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2368_2369_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2368_2369_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2368_2369_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2368_2369_add_4_1.INJECT1_1 = "NO";
    PFUMX i12294 (.BLUT(n18276), .ALUT(n14), .C0(register_addr[0]), .Z(n18278));
    LUT4 i20302_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(n26899), 
         .Z(n2650)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i20302_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut_adj_411 (.A(n79_adj_702), .B(n47), .C(n19370), .D(n26556), 
         .Z(n82)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam i1_4_lut_adj_411.init = 16'hfaea;
    RCPeripheral rc_receiver (.\register_addr[0] (register_addr[0]), .\register_addr[2] (register_addr[2]), 
            .\register_addr[1] (register_addr[1]), .\select[7] (select[7]), 
            .n176(n176), .databus_out({databus_out}), .n2(n2_adj_671), 
            .rw(rw), .databus({databus}), .\read_value[12] (read_value[12]), 
            .n1(n1_adj_667), .n28582(n28582), .\read_value[12]_adj_6 (read_value_adj_735[12]), 
            .read_value({read_value_adj_748}), .n28451(n28451), .n52(n52), 
            .n2_adj_8(n2_adj_673), .n2_adj_9(n2_adj_666), .n2_adj_10(n2_adj_662), 
            .\read_value[8]_adj_11 (read_value[8]), .n1_adj_12(n1_adj_661), 
            .\read_value[8]_adj_13 (read_value_adj_735[8]), .\read_value[9]_adj_14 (read_value[9]), 
            .n1_adj_15(n1_adj_665), .read_size({read_size}), .\read_size[0]_adj_16 (read_size_adj_789[0]), 
            .\select[1] (select[1]), .n28487(n28487), .n9(n9), .\read_size[0]_adj_17 (read_size_adj_829[0]), 
            .n28452(n28452), .n28476(n28476), .\read_size[0]_adj_18 (read_size_adj_749[0]), 
            .n10(n10), .\read_size[0]_adj_19 (read_size_adj_728[0]), .\select[2] (select[2]), 
            .n8(n8), .\read_size[2]_adj_20 (read_size_adj_789[2]), .\reg_size[2] (reg_size[2]), 
            .\read_size[2]_adj_21 (read_size_adj_829[2]), .\read_size[2]_adj_22 (read_size_adj_736[2]), 
            .\read_size[2]_adj_23 (read_size_adj_749[2]), .n28480(n28480), 
            .n4(n4_adj_652), .\read_value[0]_adj_24 (read_value_adj_828[0]), 
            .n28448(n28448), .\read_value[0]_adj_25 (read_value_adj_788[0]), 
            .\read_value[0]_adj_26 (read_value[0]), .n28458(n28458), .read_value_adj_146({read_value_adj_727}), 
            .n64(n64), .n2_adj_35(n2_adj_651), .\read_value[9]_adj_36 (read_value_adj_735[9]), 
            .n2_adj_37(n2_adj_685), .\read_value[21]_adj_38 (read_value[21]), 
            .n1_adj_39(n1_adj_684), .\read_value[31]_adj_40 (read_value[31]), 
            .n1_adj_41(n1_adj_482), .\read_value[31]_adj_42 (read_value_adj_735[31]), 
            .n4_adj_43(n4_adj_670), .\read_value[7]_adj_44 (read_value_adj_828[7]), 
            .n28576(n28576), .\sendcount[1] (sendcount[1]), .n11943(n11943), 
            .n28439(n28439), .\read_value[13]_adj_45 (read_value[13]), .n1_adj_46(n1_adj_672), 
            .n4_adj_47(n4_adj_669), .\read_value[6]_adj_48 (read_value_adj_828[6]), 
            .\read_value[7]_adj_49 (read_value_adj_788[7]), .\read_value[7]_adj_50 (read_value[7]), 
            .\read_value[13]_adj_51 (read_value_adj_735[13]), .\read_value[6]_adj_52 (read_value_adj_788[6]), 
            .\read_value[6]_adj_53 (read_value[6]), .n2_adj_54(n2_adj_664), 
            .\read_value[21]_adj_55 (read_value_adj_735[21]), .\read_value[11]_adj_56 (read_value[11]), 
            .n1_adj_57(n1_adj_663), .\read_value[10]_adj_58 (read_value_adj_735[10]), 
            .n2_adj_59(n2_adj_650), .\read_value[30]_adj_60 (read_value[30]), 
            .n1_adj_61(n1_adj_481), .n4_adj_62(n4_adj_668), .\read_value[5]_adj_63 (read_value_adj_828[5]), 
            .\read_value[5]_adj_64 (read_value_adj_788[5]), .\read_value[5]_adj_65 (read_value[5]), 
            .n30468(n30468), .\read_value[30]_adj_66 (read_value_adj_735[30]), 
            .n4_adj_67(n4_adj_658), .\read_value[4]_adj_68 (read_value_adj_828[4]), 
            .\read_value[4]_adj_69 (read_value_adj_788[4]), .\read_value[4]_adj_70 (read_value[4]), 
            .n4_adj_71(n4_adj_655), .\read_value[2]_adj_72 (read_value_adj_828[2]), 
            .\read_value[2]_adj_73 (read_value_adj_788[2]), .\read_value[2]_adj_74 (read_value[2]), 
            .\read_value[11]_adj_75 (read_value_adj_735[11]), .n2_adj_76(n2_adj_478), 
            .\read_value[28]_adj_77 (read_value[28]), .n1_adj_78(n1_adj_704), 
            .\read_value[28]_adj_79 (read_value_adj_735[28]), .n2_adj_80(n2_adj_690), 
            .\read_value[27]_adj_81 (read_value[27]), .n1_adj_82(n1_adj_696), 
            .n1_adj_83(n1_adj_656), .n2_adj_84(n2_adj_660), .\read_value[1]_adj_85 (read_value_adj_735[1]), 
            .n6(n6_adj_654), .n2_adj_86(n2_adj_681), .\read_value[20]_adj_87 (read_value[20]), 
            .n1_adj_88(n1_adj_680), .\read_value[27]_adj_89 (read_value_adj_735[27]), 
            .n2_adj_90(n2_adj_675), .\read_value[20]_adj_91 (read_value_adj_735[20]), 
            .n2_adj_92(n2_adj_677), .\read_value[14]_adj_93 (read_value[14]), 
            .n1_adj_94(n1_adj_674), .\read_value[14]_adj_95 (read_value_adj_735[14]), 
            .\read_value[19]_adj_96 (read_value[19]), .n1_adj_97(n1_adj_676), 
            .n4_adj_98(n4_adj_657), .\read_value[10]_adj_99 (read_value[10]), 
            .n1_adj_100(n1_adj_659), .\read_value[3]_adj_101 (read_value_adj_828[3]), 
            .n2_adj_102(n2_adj_484), .\read_value[19]_adj_103 (read_value_adj_735[19]), 
            .\read_value[26]_adj_104 (read_value[26]), .n1_adj_105(n1_adj_483), 
            .\read_value[3]_adj_106 (read_value_adj_788[3]), .\read_value[3]_adj_107 (read_value[3]), 
            .\read_value[26]_adj_108 (read_value_adj_735[26]), .n2_adj_109(n2_adj_480), 
            .\read_value[25]_adj_110 (read_value[25]), .n1_adj_111(n1_adj_479), 
            .n2_adj_112(n2_adj_683), .\read_value[18]_adj_113 (read_value[18]), 
            .n1_adj_114(n1_adj_682), .\read_value[25]_adj_115 (read_value_adj_735[25]), 
            .\read_value[18]_adj_116 (read_value_adj_735[18]), .n2_adj_117(n2_adj_679), 
            .\read_value[17]_adj_118 (read_value[17]), .n1_adj_119(n1_adj_678), 
            .\read_value[17]_adj_120 (read_value_adj_735[17]), .n2_adj_121(n2), 
            .\read_value[24]_adj_122 (read_value[24]), .n1_adj_123(n1), 
            .\read_value[24]_adj_124 (read_value_adj_735[24]), .\read_value[1]_adj_125 (read_value_adj_788[1]), 
            .n2_adj_126(n2_adj_689), .\read_value[16]_adj_127 (read_value[16]), 
            .n1_adj_128(n1_adj_688), .n2_adj_129(n2_adj_694), .n2_adj_130(n2_adj_700), 
            .\read_value[29]_adj_131 (read_value[29]), .n1_adj_132(n1_adj_529), 
            .\read_value[16]_adj_133 (read_value_adj_735[16]), .\read_value[29]_adj_134 (read_value_adj_735[29]), 
            .\read_value[23]_adj_135 (read_value[23]), .n1_adj_136(n1_adj_693), 
            .n2_adj_137(n2_adj_687), .\read_value[23]_adj_138 (read_value_adj_735[23]), 
            .\read_value[15]_adj_139 (read_value[15]), .n1_adj_140(n1_adj_686), 
            .n2_adj_141(n2_adj_692), .\read_value[22]_adj_142 (read_value[22]), 
            .n1_adj_143(n1_adj_691), .\read_value[15]_adj_144 (read_value_adj_735[15]), 
            .\read_value[22]_adj_145 (read_value_adj_735[22]), .debug_c_c(debug_c_c), 
            .n30470(n30470), .rc_ch8_c(rc_ch8_c), .GND_net(GND_net), .n26922(n26922), 
            .n30469(n30469), .n26942(n26942), .n12605(n12605), .n24743(n24743), 
            .n30471(n30471), .n13489(n13489), .rc_ch7_c(rc_ch7_c), .n26949(n26949), 
            .n24707(n24707), .n27040(n27040), .n13527(n13527), .rc_ch4_c(rc_ch4_c), 
            .n26947(n26947), .n24721(n24721), .n27035(n27035), .n13534(n13534), 
            .rc_ch3_c(rc_ch3_c), .n27027(n27027), .n26939(n26939), .n24755(n24755), 
            .rc_ch2_c(rc_ch2_c), .n26945(n26945), .n13535(n13535), .n24741(n24741), 
            .n27025(n27025), .n28403(n28403), .n26907(n26907), .rc_ch1_c(rc_ch1_c), 
            .n13536(n13536), .n24716(n24716), .n27023(n27023)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(621[15] 633[41])
    LUT4 i934_2_lut_3_lut (.A(n82), .B(reset_count[14]), .C(n7001), .Z(n2610)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i934_2_lut_3_lut.init = 16'hf7f7;
    PFUMX i12286 (.BLUT(n18268), .ALUT(n13), .C0(register_addr[0]), .Z(n18270));
    PFUMX i12283 (.BLUT(n18265), .ALUT(n12_adj_695), .C0(register_addr[0]), 
          .Z(n6021[3]));
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.\register_addr[1] (register_addr[1]), 
            .n24822(n24822), .debug_c_c(debug_c_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .n28477(n28477), .\read_size[0] (read_size_adj_749[0]), .n2622(n2622), 
            .n26514(n26514), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), .n12650(n12650), 
            .n579(n571_adj_766[0]), .prev_step_clk(prev_step_clk), .step_clk(step_clk), 
            .limit_latched(limit_latched_adj_531), .prev_limit_latched(prev_limit_latched_adj_532), 
            .n13363(n13363), .prev_select(prev_select_adj_567), .n28452(n28452), 
            .read_value({read_value_adj_748}), .\register_addr[0] (register_addr[0]), 
            .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), .databus({databus}), .n3539(n3539), 
            .n32(n32_adj_610), .limit_c_1(limit_c_1), .Stepper_Y_Dir_c(Stepper_Y_Dir_c), 
            .Stepper_Y_En_c(Stepper_Y_En_c), .n8273(n8273), .n611(n580_adj_767[1]), 
            .\control_reg[7] (control_reg_adj_745[7]), .n12649(n12649), 
            .n11054(n11054), .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), .\read_size[2] (read_size_adj_749[2]), 
            .n26540(n26540), .Stepper_Y_Step_c(Stepper_Y_Step_c), .n22(n22_adj_609), 
            .n28411(n28411), .n7685(n7684[7]), .n28400(n28400), .n14873(n14873), 
            .n7244(n7244), .n7278(n7278)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(573[25] 586[45])
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .read_value({read_value_adj_828}), 
            .debug_c_c(debug_c_c), .n12599(n12599), .GND_net(GND_net), 
            .n28477(n28477), .databus({databus}), .n3356(n3356), .n32(n32_adj_610), 
            .prev_step_clk(prev_step_clk), .step_clk(step_clk), .n22(n22_adj_609), 
            .VCC_net(VCC_net), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_829[0]), .n26437(n26437), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .n12795(n12795), .n579(n571_adj_766[0]), .limit_latched(limit_latched_adj_612), 
            .prev_limit_latched(prev_limit_latched_adj_613), .n12781(n12781), 
            .prev_select(prev_select_adj_648), .n28476(n28476), .n28441(n28441), 
            .n608(n580_adj_847[4]), .n610(n580_adj_847[2]), .\control_reg[7] (control_reg_adj_825[7]), 
            .n28442(n28442), .n10107(n10107), .Stepper_A_En_c(Stepper_A_En_c), 
            .Stepper_A_Dir_c(Stepper_A_Dir_c), .Stepper_A_M2_c_2(Stepper_A_M2_c_2), 
            .Stepper_A_M1_c_1(Stepper_A_M1_c_1), .\read_size[2] (read_size_adj_829[2]), 
            .n26439(n26439), .n32_adj_1(n32_adj_477), .prev_step_clk_adj_2(prev_step_clk_adj_573), 
            .step_clk_adj_3(step_clk_adj_572), .n28410(n28410), .n22_adj_4(n22), 
            .n28411(n28411), .n32_adj_5(n32), .limit_c_3(limit_c_3), .n24744(n24744), 
            .Stepper_A_Step_c(Stepper_A_Step_c), .n7703(n7702[7]), .n28399(n28399), 
            .n14876(n14876), .n7486(n7486), .n7452(n7452)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(603[25] 616[45])
    ClockDivider_U9 pwm_clk_div (.GND_net(GND_net), .n7001(n7001), .n28477(n28477), 
            .clk_255kHz(clk_255kHz), .n6966(n6966), .n26942(n26942), .n24743(n24743), 
            .n26945(n26945), .n24741(n24741), .debug_c_c(debug_c_c), .n241(n241), 
            .n26947(n26947), .n24721(n24721), .n2610(n2610), .n26949(n26949), 
            .n24707(n24707), .n26922(n26922), .n12605(n12605), .n26907(n26907), 
            .n24716(n24716), .n27027(n27027), .n13534(n13534), .n26939(n26939), 
            .n24755(n24755), .n27025(n27025), .n13535(n13535), .n27023(n27023), 
            .n13536(n13536), .n27040(n27040), .n13489(n13489), .n27035(n27035), 
            .n13527(n13527)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(518[15] 521[41])
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.debug_c_c(debug_c_c), .n28414(n28414), 
            .n28477(n28477), .databus({databus}), .n12647(n12647), .n608(n580_adj_847[4]), 
            .n610(n580_adj_847[2]), .\control_reg[7] (control_reg[7]), .n12580(n12580), 
            .n10035(n10035), .Stepper_X_En_c(Stepper_X_En_c), .Stepper_X_Dir_c(Stepper_X_Dir_c), 
            .n12583(n12583), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), .GND_net(GND_net), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\read_size[2] (read_size_adj_736[2]), 
            .n2615(n2615), .n8336(n8336), .\steps_reg[7] (steps_reg[7]), 
            .\register_addr[0] (register_addr[0]), .\read_size[0] (read_size_adj_736[0]), 
            .n28425(n28425), .Stepper_X_M0_c_0(Stepper_X_M0_c_0), .n579(n571_adj_766[0]), 
            .limit_latched(limit_latched), .prev_limit_latched(prev_limit_latched), 
            .prev_select(prev_select_adj_527), .n28480(n28480), .n3626(n3626), 
            .read_value({read_value_adj_735}), .\register_addr[1] (register_addr[1]), 
            .n19(n19), .limit_c_0(limit_c_0), .n12(n12), .VCC_net(VCC_net), 
            .Stepper_X_nFault_c(Stepper_X_nFault_c), .Stepper_X_Step_c(Stepper_X_Step_c), 
            .n24815(n24815), .n7140(n7140), .n7174(n7174), .n28401(n28401), 
            .n14714(n14714)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(558[25] 571[45])
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (\register_addr[1] , \register_addr[0] , 
            debug_c_c, n12981, n28477, databus, VCC_net, GND_net, 
            Stepper_Z_nFault_c, \read_size[0] , n13252, n233, Stepper_Z_M0_c_0, 
            n12995, n579, prev_step_clk, step_clk, limit_latched, 
            prev_limit_latched, prev_select, n28487, \read_size[2] , 
            n26489, n28438, \div_factor_reg[9] , \div_factor_reg[6] , 
            \div_factor_reg[5] , n608, n610, \control_reg[7] , n28445, 
            n10109, Stepper_Z_En_c, Stepper_Z_Dir_c, \control_reg[3] , 
            Stepper_Z_M2_c_2, Stepper_Z_M1_c_1, read_value, n3452, \steps_reg[9] , 
            \steps_reg[5] , \steps_reg[6] , \steps_reg[3] , n32, limit_c_2, 
            n24832, n6050, n18278, n18270, n79, int_step, n22, 
            n28410, \div_factor_reg[3] , n7694, n28402, n14875, n7382, 
            n7348) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[1] ;
    input \register_addr[0] ;
    input debug_c_c;
    input n12981;
    input n28477;
    input [31:0]databus;
    input VCC_net;
    input GND_net;
    input Stepper_Z_nFault_c;
    output \read_size[0] ;
    input n13252;
    input n233;
    output Stepper_Z_M0_c_0;
    input n12995;
    input n579;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    output prev_select;
    input n28487;
    output \read_size[2] ;
    input n26489;
    input n28438;
    output \div_factor_reg[9] ;
    output \div_factor_reg[6] ;
    output \div_factor_reg[5] ;
    input n608;
    input n610;
    output \control_reg[7] ;
    input n28445;
    input n10109;
    output Stepper_Z_En_c;
    output Stepper_Z_Dir_c;
    output \control_reg[3] ;
    output Stepper_Z_M2_c_2;
    output Stepper_Z_M1_c_1;
    output [31:0]read_value;
    input n3452;
    output \steps_reg[9] ;
    output \steps_reg[5] ;
    output \steps_reg[6] ;
    output \steps_reg[3] ;
    input n32;
    input limit_c_2;
    output n24832;
    input n6050;
    input n18278;
    input n18270;
    input n79;
    output int_step;
    input n22;
    input n28410;
    output \div_factor_reg[3] ;
    input n7694;
    input n28402;
    input n14875;
    output n7382;
    output n7348;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n99;
    
    wire n26808, n26809, n26810, n26820, n26821, n26822;
    wire [31:0]n100;
    
    wire fault_latched;
    wire [31:0]n3453;
    
    wire n182;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n24180;
    wire [31:0]n224;
    
    wire n24179, n24178, n24177, n24176, n24175, n26868, n26869, 
        n26870, n24174, n24173, n24172, n24171, n24170, n24169, 
        n24168, n24167, n24166, n24165;
    wire [7:0]n7693;
    wire [31:0]n5985;
    
    wire n49_adj_475, n62, n58, n50, n41_adj_476, n60, n54, n42, 
        n52, n38, n56, n46;
    wire [31:0]n6021;
    
    LUT4 i13658_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n99[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13658_4_lut.init = 16'hc088;
    LUT4 i13657_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n99[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13657_4_lut.init = 16'hc088;
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    LUT4 i13656_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n99[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13656_4_lut.init = 16'hc088;
    LUT4 i13655_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n99[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13655_4_lut.init = 16'hc088;
    PFUMX i20114 (.BLUT(n26808), .ALUT(n26809), .C0(\register_addr[1] ), 
          .Z(n26810));
    LUT4 i13654_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n99[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13654_4_lut.init = 16'hc088;
    LUT4 i13653_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n99[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13653_4_lut.init = 16'hc088;
    LUT4 i13652_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n99[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13652_4_lut.init = 16'hc088;
    LUT4 i13651_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n99[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13651_4_lut.init = 16'hc088;
    LUT4 i13650_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n99[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13650_4_lut.init = 16'hc088;
    LUT4 i13649_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n99[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13649_4_lut.init = 16'hc088;
    LUT4 i13648_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n99[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13648_4_lut.init = 16'hc088;
    LUT4 i13647_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n99[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13647_4_lut.init = 16'hc088;
    LUT4 i13646_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n99[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13646_4_lut.init = 16'hc088;
    LUT4 i13602_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n99[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13602_4_lut.init = 16'hc088;
    LUT4 i13601_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n99[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13601_4_lut.init = 16'hc088;
    LUT4 i13600_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n99[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13600_4_lut.init = 16'hc088;
    LUT4 i13599_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n99[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13599_4_lut.init = 16'hc088;
    LUT4 i13598_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n99[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13598_4_lut.init = 16'hc088;
    LUT4 i13597_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n99[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13597_4_lut.init = 16'hc088;
    LUT4 i13596_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n99[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13596_4_lut.init = 16'hc088;
    LUT4 i13595_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n99[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13595_4_lut.init = 16'hc088;
    PFUMX i20126 (.BLUT(n26820), .ALUT(n26821), .C0(\register_addr[1] ), 
          .Z(n26822));
    LUT4 i13216_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13216_4_lut.init = 16'hc088;
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3453[0]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n233), .SP(n13252), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12995), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12981), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n28487), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n26489), .SP(n13252), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3453[31]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n28438), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n28438), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n28438), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n28438), .PD(n28477), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n28438), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n28438), .PD(n28477), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n28438), .PD(n28477), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n12981), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12981), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n28445), .CD(n10109), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n28445), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n28445), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n12995), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n28445), .PD(n28477), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n12995), .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n28445), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3453[30]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3453[29]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3453[28]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3453[27]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n13252), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24180), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24179), .COUT(n24180), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24178), .COUT(n24179), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24177), .COUT(n24178), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24176), .COUT(n24177), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24175), .COUT(n24176), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    LUT4 i20124_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n26820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20124_3_lut.init = 16'hcaca;
    LUT4 i20125_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n26821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20125_3_lut.init = 16'hcaca;
    PFUMX i20174 (.BLUT(n26868), .ALUT(n26869), .C0(\register_addr[0] ), 
          .Z(n26870));
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24174), .COUT(n24175), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24173), .COUT(n24174), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24172), .COUT(n24173), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24171), .COUT(n24172), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    LUT4 mux_1471_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3452), .Z(n3453[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i1_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24170), .COUT(n24171), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24169), .COUT(n24170), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24168), .COUT(n24169), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24167), .COUT(n24168), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24166), .COUT(n24167), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24165), .COUT(n24166), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n24165), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i13215_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7693[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13215_2_lut.init = 16'h2222;
    LUT4 mux_1781_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5985[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1781_i5_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i26 (.D(n3453[26]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    LUT4 mux_1781_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5985[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1781_i8_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i25 (.D(n3453[25]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3453[24]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3453[23]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3453[22]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3453[21]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3453[20]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3453[19]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3453[18]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3453[17]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3453[16]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3453[15]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3453[14]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3453[13]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3453[12]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3453[11]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3453[10]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3453[9]), .CK(debug_c_c), .CD(n28477), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3453[8]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3453[7]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3453[6]), .CK(debug_c_c), .CD(n28477), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3453[5]), .CK(debug_c_c), .CD(n28477), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3453[4]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3453[3]), .CK(debug_c_c), .CD(n28477), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3453[2]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3453[1]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i13659_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n99[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13659_4_lut.init = 16'hc088;
    LUT4 i20172_3_lut (.A(Stepper_Z_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n26868)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20172_3_lut.init = 16'hcaca;
    LUT4 i20173_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n26869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20173_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49_adj_475), .B(n62), .C(n58), .D(n50), .Z(n24832)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49_adj_475)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41_adj_476), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41_adj_476)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 mux_1471_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3452), 
         .Z(n3453[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i32_3_lut.init = 16'hcaca;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    FD1P3IX read_value__i1 (.D(n26822), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n26870), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6050), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6021[4]), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18278), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n18270), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6021[7]), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n99[8]), .SP(n13252), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n79), .SP(n13252), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n99[10]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n99[11]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n99[12]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n99[13]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n99[14]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n99[15]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n99[16]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n99[17]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n99[18]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n99[19]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n99[20]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n99[21]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n99[22]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n99[23]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n99[24]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n99[25]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n99[26]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n99[27]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n99[28]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n99[29]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n99[30]), .SP(n13252), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n28410), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n26810), .SP(n13252), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    PFUMX mux_1785_i5 (.BLUT(n7693[4]), .ALUT(n5985[4]), .C0(\register_addr[1] ), 
          .Z(n6021[4]));
    PFUMX mux_1785_i8 (.BLUT(n7694), .ALUT(n5985[7]), .C0(\register_addr[1] ), 
          .Z(n6021[7]));
    LUT4 mux_1471_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3452), 
         .Z(n3453[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3452), 
         .Z(n3453[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3452), 
         .Z(n3453[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3452), 
         .Z(n3453[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3452), 
         .Z(n3453[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3452), 
         .Z(n3453[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3452), 
         .Z(n3453[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3452), 
         .Z(n3453[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3452), 
         .Z(n3453[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3452), 
         .Z(n3453[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3452), 
         .Z(n3453[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3452), 
         .Z(n3453[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3452), 
         .Z(n3453[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3452), 
         .Z(n3453[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3452), 
         .Z(n3453[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3452), 
         .Z(n3453[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i12_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    LUT4 mux_1471_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3452), 
         .Z(n3453[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3452), .Z(n3453[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3452), .Z(n3453[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3452), .Z(n3453[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3452), .Z(n3453[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3452), .Z(n3453[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3452), .Z(n3453[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3452), .Z(n3453[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3452), .Z(n3453[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3452), .Z(n3453[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3452), 
         .Z(n3453[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3452), 
         .Z(n3453[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3452), 
         .Z(n3453[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1471_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3452), 
         .Z(n3453[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1471_i28_3_lut.init = 16'hcaca;
    LUT4 i20112_3_lut (.A(Stepper_Z_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n26808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20112_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    LUT4 i20113_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n26809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20113_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12981), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    ClockDivider step_clk_gen (.GND_net(GND_net), .div_factor_reg({div_factor_reg[31:10], 
            \div_factor_reg[9] , div_factor_reg[8:7], \div_factor_reg[6] , 
            \div_factor_reg[5] , div_factor_reg[4], \div_factor_reg[3] , 
            div_factor_reg[2:0]}), .step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n28477(n28477), .n28402(n28402), .n14875(n14875), .n7382(n7382), 
            .n7348(n7348)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (GND_net, div_factor_reg, step_clk, debug_c_c, n28477, 
            n28402, n14875, n7382, n7348) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [31:0]div_factor_reg;
    output step_clk;
    input debug_c_c;
    input n28477;
    input n28402;
    input n14875;
    output n7382;
    output n7348;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n23845, n7313;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n23908, n23907, n23906, n23905, n23904, n23903, n23902, 
        n23901, n23900, n23899, n23898, n23897, n23896, n23895, 
        n23860, n23894, n23893, n24116;
    wire [31:0]n40;
    
    wire n24115, n24114, n24113, n24112, n24111, n24110, n24109, 
        n23892, n24108, n24107, n23859, n23858, n23891, n24106, 
        n24105, n23857, n23890, n24104, n24103, n23889, n24102, 
        n23856, n23888, n24101, n23887, n23855, n23886, n23854, 
        n24248, n23885, n24247, n24246, n24245, n24244, n23884, 
        n24243, n24242, n24241, n23853, n24240, n24239, n24238, 
        n24237, n23883, n23852, n24236, n24235, n24234, n24233, 
        n23882, n23851, n23850, n23881, n23849, n23880, n23848, 
        n23847, n23879, n23878, n23877, n23846;
    
    CCU2D sub_1879_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n23845));
    defparam sub_1879_add_2_1.INIT0 = 16'h0000;
    defparam sub_1879_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1879_add_2_1.INJECT1_0 = "NO";
    defparam sub_1879_add_2_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7313), .CK(debug_c_c), .CD(n28477), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2374__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    CCU2D sub_1876_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23908), .S1(n7313));
    defparam sub_1876_add_2_33.INIT0 = 16'h5555;
    defparam sub_1876_add_2_33.INIT1 = 16'h0000;
    defparam sub_1876_add_2_33.INJECT1_0 = "NO";
    defparam sub_1876_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23907), .COUT(n23908));
    defparam sub_1876_add_2_31.INIT0 = 16'h5999;
    defparam sub_1876_add_2_31.INIT1 = 16'h5999;
    defparam sub_1876_add_2_31.INJECT1_0 = "NO";
    defparam sub_1876_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28402), .PD(n14875), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_1876_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23906), .COUT(n23907));
    defparam sub_1876_add_2_29.INIT0 = 16'h5999;
    defparam sub_1876_add_2_29.INIT1 = 16'h5999;
    defparam sub_1876_add_2_29.INJECT1_0 = "NO";
    defparam sub_1876_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23905), .COUT(n23906));
    defparam sub_1876_add_2_27.INIT0 = 16'h5999;
    defparam sub_1876_add_2_27.INIT1 = 16'h5999;
    defparam sub_1876_add_2_27.INJECT1_0 = "NO";
    defparam sub_1876_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23904), .COUT(n23905));
    defparam sub_1876_add_2_25.INIT0 = 16'h5999;
    defparam sub_1876_add_2_25.INIT1 = 16'h5999;
    defparam sub_1876_add_2_25.INJECT1_0 = "NO";
    defparam sub_1876_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23903), .COUT(n23904));
    defparam sub_1876_add_2_23.INIT0 = 16'h5999;
    defparam sub_1876_add_2_23.INIT1 = 16'h5999;
    defparam sub_1876_add_2_23.INJECT1_0 = "NO";
    defparam sub_1876_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23902), .COUT(n23903));
    defparam sub_1876_add_2_21.INIT0 = 16'h5999;
    defparam sub_1876_add_2_21.INIT1 = 16'h5999;
    defparam sub_1876_add_2_21.INJECT1_0 = "NO";
    defparam sub_1876_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23901), .COUT(n23902));
    defparam sub_1876_add_2_19.INIT0 = 16'h5999;
    defparam sub_1876_add_2_19.INIT1 = 16'h5999;
    defparam sub_1876_add_2_19.INJECT1_0 = "NO";
    defparam sub_1876_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23900), .COUT(n23901));
    defparam sub_1876_add_2_17.INIT0 = 16'h5999;
    defparam sub_1876_add_2_17.INIT1 = 16'h5999;
    defparam sub_1876_add_2_17.INJECT1_0 = "NO";
    defparam sub_1876_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23899), .COUT(n23900));
    defparam sub_1876_add_2_15.INIT0 = 16'h5999;
    defparam sub_1876_add_2_15.INIT1 = 16'h5999;
    defparam sub_1876_add_2_15.INJECT1_0 = "NO";
    defparam sub_1876_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23898), .COUT(n23899));
    defparam sub_1876_add_2_13.INIT0 = 16'h5999;
    defparam sub_1876_add_2_13.INIT1 = 16'h5999;
    defparam sub_1876_add_2_13.INJECT1_0 = "NO";
    defparam sub_1876_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23897), .COUT(n23898));
    defparam sub_1876_add_2_11.INIT0 = 16'h5999;
    defparam sub_1876_add_2_11.INIT1 = 16'h5999;
    defparam sub_1876_add_2_11.INJECT1_0 = "NO";
    defparam sub_1876_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23896), .COUT(n23897));
    defparam sub_1876_add_2_9.INIT0 = 16'h5999;
    defparam sub_1876_add_2_9.INIT1 = 16'h5999;
    defparam sub_1876_add_2_9.INJECT1_0 = "NO";
    defparam sub_1876_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23895), .COUT(n23896));
    defparam sub_1876_add_2_7.INIT0 = 16'h5999;
    defparam sub_1876_add_2_7.INIT1 = 16'h5999;
    defparam sub_1876_add_2_7.INJECT1_0 = "NO";
    defparam sub_1876_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23860), .S1(n7382));
    defparam sub_1879_add_2_33.INIT0 = 16'hf555;
    defparam sub_1879_add_2_33.INIT1 = 16'h0000;
    defparam sub_1879_add_2_33.INJECT1_0 = "NO";
    defparam sub_1879_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23894), .COUT(n23895));
    defparam sub_1876_add_2_5.INIT0 = 16'h5999;
    defparam sub_1876_add_2_5.INIT1 = 16'h5999;
    defparam sub_1876_add_2_5.INJECT1_0 = "NO";
    defparam sub_1876_add_2_5.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28402), .CD(n14875), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1S3IX count_2374__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i1.GSR = "ENABLED";
    FD1S3IX count_2374__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i2.GSR = "ENABLED";
    FD1S3IX count_2374__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i3.GSR = "ENABLED";
    FD1S3IX count_2374__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i4.GSR = "ENABLED";
    FD1S3IX count_2374__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i5.GSR = "ENABLED";
    FD1S3IX count_2374__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i6.GSR = "ENABLED";
    FD1S3IX count_2374__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i7.GSR = "ENABLED";
    FD1S3IX count_2374__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i8.GSR = "ENABLED";
    FD1S3IX count_2374__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i9.GSR = "ENABLED";
    FD1S3IX count_2374__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i10.GSR = "ENABLED";
    FD1S3IX count_2374__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i11.GSR = "ENABLED";
    FD1S3IX count_2374__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i12.GSR = "ENABLED";
    FD1S3IX count_2374__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i13.GSR = "ENABLED";
    FD1S3IX count_2374__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i14.GSR = "ENABLED";
    FD1S3IX count_2374__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i15.GSR = "ENABLED";
    FD1S3IX count_2374__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i16.GSR = "ENABLED";
    FD1S3IX count_2374__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i17.GSR = "ENABLED";
    FD1S3IX count_2374__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i18.GSR = "ENABLED";
    FD1S3IX count_2374__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i19.GSR = "ENABLED";
    FD1S3IX count_2374__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i20.GSR = "ENABLED";
    FD1S3IX count_2374__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i21.GSR = "ENABLED";
    FD1S3IX count_2374__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i22.GSR = "ENABLED";
    FD1S3IX count_2374__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i23.GSR = "ENABLED";
    FD1S3IX count_2374__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i24.GSR = "ENABLED";
    FD1S3IX count_2374__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i25.GSR = "ENABLED";
    FD1S3IX count_2374__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i26.GSR = "ENABLED";
    FD1S3IX count_2374__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i27.GSR = "ENABLED";
    FD1S3IX count_2374__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i28.GSR = "ENABLED";
    FD1S3IX count_2374__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i29.GSR = "ENABLED";
    FD1S3IX count_2374__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i30.GSR = "ENABLED";
    FD1S3IX count_2374__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28402), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374__i31.GSR = "ENABLED";
    CCU2D sub_1876_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23893), .COUT(n23894));
    defparam sub_1876_add_2_3.INIT0 = 16'h5999;
    defparam sub_1876_add_2_3.INIT1 = 16'h5999;
    defparam sub_1876_add_2_3.INJECT1_0 = "NO";
    defparam sub_1876_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1876_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n23893));
    defparam sub_1876_add_2_1.INIT0 = 16'h0000;
    defparam sub_1876_add_2_1.INIT1 = 16'h5999;
    defparam sub_1876_add_2_1.INJECT1_0 = "NO";
    defparam sub_1876_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24116), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24115), .COUT(n24116), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24114), .COUT(n24115), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24113), .COUT(n24114), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24112), .COUT(n24113), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24111), .COUT(n24112), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24110), .COUT(n24111), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24109), .COUT(n24110), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23892), .S1(n7348));
    defparam sub_1878_add_2_33.INIT0 = 16'h5999;
    defparam sub_1878_add_2_33.INIT1 = 16'h0000;
    defparam sub_1878_add_2_33.INJECT1_0 = "NO";
    defparam sub_1878_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24108), .COUT(n24109), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24107), .COUT(n24108), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23859), .COUT(n23860));
    defparam sub_1879_add_2_31.INIT0 = 16'hf555;
    defparam sub_1879_add_2_31.INIT1 = 16'hf555;
    defparam sub_1879_add_2_31.INJECT1_0 = "NO";
    defparam sub_1879_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23858), .COUT(n23859));
    defparam sub_1879_add_2_29.INIT0 = 16'hf555;
    defparam sub_1879_add_2_29.INIT1 = 16'hf555;
    defparam sub_1879_add_2_29.INJECT1_0 = "NO";
    defparam sub_1879_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23891), .COUT(n23892));
    defparam sub_1878_add_2_31.INIT0 = 16'h5999;
    defparam sub_1878_add_2_31.INIT1 = 16'h5999;
    defparam sub_1878_add_2_31.INJECT1_0 = "NO";
    defparam sub_1878_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24106), .COUT(n24107), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24105), .COUT(n24106), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23857), .COUT(n23858));
    defparam sub_1879_add_2_27.INIT0 = 16'hf555;
    defparam sub_1879_add_2_27.INIT1 = 16'hf555;
    defparam sub_1879_add_2_27.INJECT1_0 = "NO";
    defparam sub_1879_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23890), .COUT(n23891));
    defparam sub_1878_add_2_29.INIT0 = 16'h5999;
    defparam sub_1878_add_2_29.INIT1 = 16'h5999;
    defparam sub_1878_add_2_29.INJECT1_0 = "NO";
    defparam sub_1878_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24104), .COUT(n24105), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24103), .COUT(n24104), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23889), .COUT(n23890));
    defparam sub_1878_add_2_27.INIT0 = 16'h5999;
    defparam sub_1878_add_2_27.INIT1 = 16'h5999;
    defparam sub_1878_add_2_27.INJECT1_0 = "NO";
    defparam sub_1878_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24102), .COUT(n24103), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23856), .COUT(n23857));
    defparam sub_1879_add_2_25.INIT0 = 16'hf555;
    defparam sub_1879_add_2_25.INIT1 = 16'hf555;
    defparam sub_1879_add_2_25.INJECT1_0 = "NO";
    defparam sub_1879_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23888), .COUT(n23889));
    defparam sub_1878_add_2_25.INIT0 = 16'h5999;
    defparam sub_1878_add_2_25.INIT1 = 16'h5999;
    defparam sub_1878_add_2_25.INJECT1_0 = "NO";
    defparam sub_1878_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24101), .COUT(n24102), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23887), .COUT(n23888));
    defparam sub_1878_add_2_23.INIT0 = 16'h5999;
    defparam sub_1878_add_2_23.INIT1 = 16'h5999;
    defparam sub_1878_add_2_23.INJECT1_0 = "NO";
    defparam sub_1878_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23855), .COUT(n23856));
    defparam sub_1879_add_2_23.INIT0 = 16'hf555;
    defparam sub_1879_add_2_23.INIT1 = 16'hf555;
    defparam sub_1879_add_2_23.INJECT1_0 = "NO";
    defparam sub_1879_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23886), .COUT(n23887));
    defparam sub_1878_add_2_21.INIT0 = 16'h5999;
    defparam sub_1878_add_2_21.INIT1 = 16'h5999;
    defparam sub_1878_add_2_21.INJECT1_0 = "NO";
    defparam sub_1878_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23854), .COUT(n23855));
    defparam sub_1879_add_2_21.INIT0 = 16'hf555;
    defparam sub_1879_add_2_21.INIT1 = 16'hf555;
    defparam sub_1879_add_2_21.INJECT1_0 = "NO";
    defparam sub_1879_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24248), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_33.INIT1 = 16'h0000;
    defparam count_2374_add_4_33.INJECT1_0 = "NO";
    defparam count_2374_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24101), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23885), .COUT(n23886));
    defparam sub_1878_add_2_19.INIT0 = 16'h5999;
    defparam sub_1878_add_2_19.INIT1 = 16'h5999;
    defparam sub_1878_add_2_19.INJECT1_0 = "NO";
    defparam sub_1878_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24247), .COUT(n24248), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_31.INJECT1_0 = "NO";
    defparam count_2374_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24246), .COUT(n24247), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_29.INJECT1_0 = "NO";
    defparam count_2374_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24245), .COUT(n24246), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_27.INJECT1_0 = "NO";
    defparam count_2374_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24244), .COUT(n24245), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_25.INJECT1_0 = "NO";
    defparam count_2374_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23884), .COUT(n23885));
    defparam sub_1878_add_2_17.INIT0 = 16'h5999;
    defparam sub_1878_add_2_17.INIT1 = 16'h5999;
    defparam sub_1878_add_2_17.INJECT1_0 = "NO";
    defparam sub_1878_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24243), .COUT(n24244), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_23.INJECT1_0 = "NO";
    defparam count_2374_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24242), .COUT(n24243), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_21.INJECT1_0 = "NO";
    defparam count_2374_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24241), .COUT(n24242), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_19.INJECT1_0 = "NO";
    defparam count_2374_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23853), .COUT(n23854));
    defparam sub_1879_add_2_19.INIT0 = 16'hf555;
    defparam sub_1879_add_2_19.INIT1 = 16'hf555;
    defparam sub_1879_add_2_19.INJECT1_0 = "NO";
    defparam sub_1879_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24240), .COUT(n24241), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_17.INJECT1_0 = "NO";
    defparam count_2374_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24239), .COUT(n24240), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_15.INJECT1_0 = "NO";
    defparam count_2374_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24238), .COUT(n24239), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_13.INJECT1_0 = "NO";
    defparam count_2374_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24237), .COUT(n24238), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_11.INJECT1_0 = "NO";
    defparam count_2374_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23883), .COUT(n23884));
    defparam sub_1878_add_2_15.INIT0 = 16'h5999;
    defparam sub_1878_add_2_15.INIT1 = 16'h5999;
    defparam sub_1878_add_2_15.INJECT1_0 = "NO";
    defparam sub_1878_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23852), .COUT(n23853));
    defparam sub_1879_add_2_17.INIT0 = 16'hf555;
    defparam sub_1879_add_2_17.INIT1 = 16'hf555;
    defparam sub_1879_add_2_17.INJECT1_0 = "NO";
    defparam sub_1879_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24236), .COUT(n24237), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_9.INJECT1_0 = "NO";
    defparam count_2374_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24235), .COUT(n24236), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_7.INJECT1_0 = "NO";
    defparam count_2374_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24234), .COUT(n24235), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_5.INJECT1_0 = "NO";
    defparam count_2374_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24233), .COUT(n24234), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2374_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2374_add_4_3.INJECT1_0 = "NO";
    defparam count_2374_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2374_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24233), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2374_add_4_1.INIT0 = 16'hF000;
    defparam count_2374_add_4_1.INIT1 = 16'h0555;
    defparam count_2374_add_4_1.INJECT1_0 = "NO";
    defparam count_2374_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23882), .COUT(n23883));
    defparam sub_1878_add_2_13.INIT0 = 16'h5999;
    defparam sub_1878_add_2_13.INIT1 = 16'h5999;
    defparam sub_1878_add_2_13.INJECT1_0 = "NO";
    defparam sub_1878_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23851), .COUT(n23852));
    defparam sub_1879_add_2_15.INIT0 = 16'hf555;
    defparam sub_1879_add_2_15.INIT1 = 16'hf555;
    defparam sub_1879_add_2_15.INJECT1_0 = "NO";
    defparam sub_1879_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23850), .COUT(n23851));
    defparam sub_1879_add_2_13.INIT0 = 16'hf555;
    defparam sub_1879_add_2_13.INIT1 = 16'hf555;
    defparam sub_1879_add_2_13.INJECT1_0 = "NO";
    defparam sub_1879_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23881), .COUT(n23882));
    defparam sub_1878_add_2_11.INIT0 = 16'h5999;
    defparam sub_1878_add_2_11.INIT1 = 16'h5999;
    defparam sub_1878_add_2_11.INJECT1_0 = "NO";
    defparam sub_1878_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23849), .COUT(n23850));
    defparam sub_1879_add_2_11.INIT0 = 16'hf555;
    defparam sub_1879_add_2_11.INIT1 = 16'hf555;
    defparam sub_1879_add_2_11.INJECT1_0 = "NO";
    defparam sub_1879_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23880), .COUT(n23881));
    defparam sub_1878_add_2_9.INIT0 = 16'h5999;
    defparam sub_1878_add_2_9.INIT1 = 16'h5999;
    defparam sub_1878_add_2_9.INJECT1_0 = "NO";
    defparam sub_1878_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23848), .COUT(n23849));
    defparam sub_1879_add_2_9.INIT0 = 16'hf555;
    defparam sub_1879_add_2_9.INIT1 = 16'hf555;
    defparam sub_1879_add_2_9.INJECT1_0 = "NO";
    defparam sub_1879_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23847), .COUT(n23848));
    defparam sub_1879_add_2_7.INIT0 = 16'hf555;
    defparam sub_1879_add_2_7.INIT1 = 16'hf555;
    defparam sub_1879_add_2_7.INJECT1_0 = "NO";
    defparam sub_1879_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23879), .COUT(n23880));
    defparam sub_1878_add_2_7.INIT0 = 16'h5999;
    defparam sub_1878_add_2_7.INIT1 = 16'h5999;
    defparam sub_1878_add_2_7.INJECT1_0 = "NO";
    defparam sub_1878_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23878), .COUT(n23879));
    defparam sub_1878_add_2_5.INIT0 = 16'h5999;
    defparam sub_1878_add_2_5.INIT1 = 16'h5999;
    defparam sub_1878_add_2_5.INJECT1_0 = "NO";
    defparam sub_1878_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23877), .COUT(n23878));
    defparam sub_1878_add_2_3.INIT0 = 16'h5999;
    defparam sub_1878_add_2_3.INIT1 = 16'h5999;
    defparam sub_1878_add_2_3.INJECT1_0 = "NO";
    defparam sub_1878_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1878_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n23877));
    defparam sub_1878_add_2_1.INIT0 = 16'h0000;
    defparam sub_1878_add_2_1.INIT1 = 16'h5999;
    defparam sub_1878_add_2_1.INJECT1_0 = "NO";
    defparam sub_1878_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23846), .COUT(n23847));
    defparam sub_1879_add_2_5.INIT0 = 16'hf555;
    defparam sub_1879_add_2_5.INIT1 = 16'hf555;
    defparam sub_1879_add_2_5.INJECT1_0 = "NO";
    defparam sub_1879_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1879_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23845), .COUT(n23846));
    defparam sub_1879_add_2_3.INIT0 = 16'hf555;
    defparam sub_1879_add_2_3.INIT1 = 16'hf555;
    defparam sub_1879_add_2_3.INJECT1_0 = "NO";
    defparam sub_1879_add_2_3.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (debug_c_c, n8430, n28477, read_size, 
            n12585, n19316, prev_clk_1Hz, clk_1Hz, prev_select, \select[1] , 
            xbee_pause_c, n28537, \register[1][1] , n28504, \control_reg[7] , 
            n24822, n32, \control_reg[7]_adj_238 , n24815, n19, \register[0][7] , 
            n28508, n19865, n28505, \register[1][7] , n28506, n19338, 
            \register[0][4] , n17481, \control_reg[7]_adj_239 , n24744, 
            n32_adj_240, \register[2][31] , \register[2][30] , \register[2][29] , 
            \register[2][28] , \register[2][27] , \register[2][26] , \register[2][25] , 
            \register[2][24] , \register[2][23] , \register[2][22] , \register[2][21] , 
            \register[2][20] , \register[2][19] , \register[2][18] , \register[2][17] , 
            \register[2][16] , \register[2][15] , \register[2][14] , \register[2][13] , 
            \register[2][12] , \register[2][11] , \register[2][10] , \register[2][9] , 
            \register[2][8] , \register[2][7] , \register[2][6] , \register[2][5] , 
            \register[2][4] , \control_reg[7]_adj_241 , n24832, n32_adj_242, 
            signal_light_c, \register_addr[1] , \register_addr[0] , n27504, 
            n27502, n11, n28431, rw, n15, n28582, n6, \read_value[2] , 
            n27505, n27503, \read_value[3] , n8472, \read_value[4] , 
            n26100, \read_value[5] , n26096, \read_value[6] , n26088, 
            \read_value[7] , n26090, \read_value[8] , n26076, \read_value[9] , 
            n26077, \read_value[10] , n26081, \read_value[11] , n26083, 
            \read_value[12] , n26098, \read_value[13] , n26085, \read_value[14] , 
            n26079, \read_value[15] , n26087, \read_value[16] , n26084, 
            \read_value[17] , n26094, \read_value[18] , n26095, \read_value[19] , 
            n26093, \read_value[20] , n26091, \read_value[21] , n26092, 
            \read_value[22] , n26080, \read_value[23] , n26086, \read_value[24] , 
            n26078, \read_value[25] , n26082, \read_value[26] , n26089, 
            \read_value[27] , n26102, \read_value[28] , n26097, \read_value[29] , 
            n26099, \read_value[30] , n26103, \read_value[31] , n26101, 
            \databus[1] , GND_net, n26425, n62, n14798, n15_adj_243, 
            \read_value[0] , n4, n2650, n26899) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n8430;
    input n28477;
    output [2:0]read_size;
    input n12585;
    input n19316;
    output prev_clk_1Hz;
    output clk_1Hz;
    output prev_select;
    input \select[1] ;
    input xbee_pause_c;
    output n28537;
    input \register[1][1] ;
    output n28504;
    input \control_reg[7] ;
    input n24822;
    output n32;
    input \control_reg[7]_adj_238 ;
    input n24815;
    output n19;
    input \register[0][7] ;
    output n28508;
    input n19865;
    output n28505;
    input \register[1][7] ;
    output n28506;
    output n19338;
    input \register[0][4] ;
    output n17481;
    input \control_reg[7]_adj_239 ;
    input n24744;
    output n32_adj_240;
    output \register[2][31] ;
    output \register[2][30] ;
    output \register[2][29] ;
    output \register[2][28] ;
    output \register[2][27] ;
    output \register[2][26] ;
    output \register[2][25] ;
    output \register[2][24] ;
    output \register[2][23] ;
    output \register[2][22] ;
    output \register[2][21] ;
    output \register[2][20] ;
    output \register[2][19] ;
    output \register[2][18] ;
    output \register[2][17] ;
    output \register[2][16] ;
    output \register[2][15] ;
    output \register[2][14] ;
    output \register[2][13] ;
    output \register[2][12] ;
    output \register[2][11] ;
    output \register[2][10] ;
    output \register[2][9] ;
    output \register[2][8] ;
    output \register[2][7] ;
    output \register[2][6] ;
    output \register[2][5] ;
    output \register[2][4] ;
    input \control_reg[7]_adj_241 ;
    input n24832;
    output n32_adj_242;
    output signal_light_c;
    input \register_addr[1] ;
    input \register_addr[0] ;
    output n27504;
    output n27502;
    output n11;
    input n28431;
    input rw;
    input n15;
    output n28582;
    output n6;
    output \read_value[2] ;
    input n27505;
    input n27503;
    output \read_value[3] ;
    input n8472;
    output \read_value[4] ;
    input n26100;
    output \read_value[5] ;
    input n26096;
    output \read_value[6] ;
    input n26088;
    output \read_value[7] ;
    input n26090;
    output \read_value[8] ;
    input n26076;
    output \read_value[9] ;
    input n26077;
    output \read_value[10] ;
    input n26081;
    output \read_value[11] ;
    input n26083;
    output \read_value[12] ;
    input n26098;
    output \read_value[13] ;
    input n26085;
    output \read_value[14] ;
    input n26079;
    output \read_value[15] ;
    input n26087;
    output \read_value[16] ;
    input n26084;
    output \read_value[17] ;
    input n26094;
    output \read_value[18] ;
    input n26095;
    output \read_value[19] ;
    input n26093;
    output \read_value[20] ;
    input n26091;
    output \read_value[21] ;
    input n26092;
    output \read_value[22] ;
    input n26080;
    output \read_value[23] ;
    input n26086;
    output \read_value[24] ;
    input n26078;
    output \read_value[25] ;
    input n26082;
    output \read_value[26] ;
    input n26089;
    output \read_value[27] ;
    input n26102;
    output \read_value[28] ;
    input n26097;
    output \read_value[29] ;
    input n26099;
    output \read_value[30] ;
    input n26103;
    output \read_value[31] ;
    input n26101;
    input \databus[1] ;
    input GND_net;
    input n26425;
    input n62;
    input n14798;
    input n15_adj_243;
    output \read_value[0] ;
    input n4;
    input n2650;
    output n26899;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    wire [31:0]n100;
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n178, force_pause, n10231, n26772;
    wire [31:0]n6739;
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    
    wire n25341, n24020, n24019, n24018, n24017, n24016, n24015, 
        n24014, n24013, n24012, n24011, n24010, n24009, n24008, 
        n24007, n24006, n24005;
    
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n19316), .SP(n12585), .CK(debug_c_c), 
            .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_149 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_clk_1Hz_149.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_150 (.D(n178), .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam xbee_pause_latched_150.GSR = "ENABLED";
    FD1S3AX prev_select_148 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_select_148.GSR = "ENABLED";
    LUT4 i114_1_lut (.A(xbee_pause_c), .Z(n178)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(54[26:39])
    defparam i114_1_lut.init = 16'h5555;
    LUT4 i112_2_lut_rep_416 (.A(\register[0] [2]), .B(force_pause), .Z(n28537)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i112_2_lut_rep_416.init = 16'heeee;
    LUT4 i13136_2_lut_rep_383_3_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(\register[1][1] ), .Z(n28504)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i13136_2_lut_rep_383_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(\control_reg[7] ), 
         .D(n24822), .Z(n32)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_398 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_238 ), .D(n24815), .Z(n19)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_398.init = 16'h1000;
    LUT4 i13130_2_lut_rep_387_3_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(\register[0][7] ), .Z(n28508)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i13130_2_lut_rep_387_3_lut.init = 16'h1010;
    LUT4 i13884_2_lut_rep_384_4_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(n19865), .D(\register[1][1] ), .Z(n28505)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i13884_2_lut_rep_384_4_lut.init = 16'hf0e0;
    LUT4 i13132_2_lut_rep_385_3_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(\register[1][7] ), .Z(n28506)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i13132_2_lut_rep_385_3_lut.init = 16'h1010;
    LUT4 i20369_2_lut_2_lut_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(n19865), .D(\register[1][1] ), .Z(n19338)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i20369_2_lut_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i1_3_lut_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(\register[0][4] ), 
         .D(\register[0][7] ), .Z(n17481)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_399 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_239 ), .D(n24744), .Z(n32_adj_240)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_399.init = 16'h1000;
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][31] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][30] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][29] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][28] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][27] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][26] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][25] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][23] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][22] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][21] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][19] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][18] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][17] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n8430), .CD(n28477), 
            .CK(debug_c_c), .Q(\register[2][10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2][9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2][8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2][7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2][6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2][5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    LUT4 i2_3_lut_4_lut_adj_400 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_241 ), .D(n24832), .Z(n32_adj_242)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_400.init = 16'h1000;
    LUT4 i13101_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(clk_1Hz), 
         .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i13101_2_lut_3_lut.init = 16'hfefe;
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n8430), .CD(n28477), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    LUT4 i4231_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(\register_addr[1] ), 
         .D(\register[2] [0]), .Z(n10231)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i4231_3_lut_4_lut.init = 16'hfe0e;
    LUT4 register_addr_0__bdd_4_lut (.A(\register_addr[0] ), .B(\register[0] [2]), 
         .C(\register_addr[1] ), .D(\register[2] [2]), .Z(n27504)) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam register_addr_0__bdd_4_lut.init = 16'h5e0e;
    LUT4 register_addr_0__bdd_4_lut_20572 (.A(\register_addr[0] ), .B(force_pause), 
         .C(\register_addr[1] ), .D(\register[2] [1]), .Z(n27502)) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam register_addr_0__bdd_4_lut_20572.init = 16'h5e0e;
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n11)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i20078_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n28431), .C(prev_select), 
         .D(rw), .Z(n26772)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20078_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i13064_4_lut (.A(n28431), .B(n15), .C(n10231), .D(\register_addr[0] ), 
         .Z(n6739[0])) /* synthesis lut_function=(!(A (B)+!A (B ((D)+!C)))) */ ;
    defparam i13064_4_lut.init = 16'h3373;
    LUT4 i14_2_lut_rep_461 (.A(\select[1] ), .B(rw), .Z(n28582)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam i14_2_lut_rep_461.init = 16'h8888;
    LUT4 Select_3960_i6_2_lut_3_lut (.A(\select[1] ), .B(rw), .C(read_value[1]), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam Select_3960_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_4_lut (.A(\select[1] ), .B(n28477), .C(n26772), .D(\register_addr[0] ), 
         .Z(n25341)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccce;
    FD1P3AX read_value__i2 (.D(n27505), .SP(n12585), .CK(debug_c_c), .Q(\read_value[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3AX read_value__i1 (.D(n27503), .SP(n12585), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6739[3]), .SP(n12585), .CD(n8472), .CK(debug_c_c), 
            .Q(\read_value[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n26100), .SP(n12585), .CK(debug_c_c), .Q(\read_value[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n26096), .SP(n12585), .CK(debug_c_c), .Q(\read_value[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n26088), .SP(n12585), .CK(debug_c_c), .Q(\read_value[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n26090), .SP(n12585), .CK(debug_c_c), .Q(\read_value[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n26076), .SP(n12585), .CK(debug_c_c), .Q(\read_value[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n26077), .SP(n12585), .CK(debug_c_c), .Q(\read_value[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n26081), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n26083), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n26098), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n26085), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n26079), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n26087), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n26084), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n26094), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[17] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n26095), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[18] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n26093), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[19] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n26091), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n26092), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[21] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n26080), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[22] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n26086), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[23] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n26078), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n26082), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[25] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n26089), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[26] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n26102), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[27] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n26097), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[28] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n26099), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[29] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n26103), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[30] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n26101), .SP(n12585), .CK(debug_c_c), 
            .Q(\read_value[31] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX force_pause_151 (.D(\databus[1] ), .SP(n25341), .CD(n28477), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam force_pause_151.GSR = "ENABLED";
    CCU2D add_134_33 (.A0(\register[2][31] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24020), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_33.INIT0 = 16'h5aaa;
    defparam add_134_33.INIT1 = 16'h0000;
    defparam add_134_33.INJECT1_0 = "NO";
    defparam add_134_33.INJECT1_1 = "NO";
    CCU2D add_134_31 (.A0(\register[2][29] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][30] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24019), .COUT(n24020), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_31.INIT0 = 16'h5aaa;
    defparam add_134_31.INIT1 = 16'h5aaa;
    defparam add_134_31.INJECT1_0 = "NO";
    defparam add_134_31.INJECT1_1 = "NO";
    CCU2D add_134_29 (.A0(\register[2][27] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][28] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24018), .COUT(n24019), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_29.INIT0 = 16'h5aaa;
    defparam add_134_29.INIT1 = 16'h5aaa;
    defparam add_134_29.INJECT1_0 = "NO";
    defparam add_134_29.INJECT1_1 = "NO";
    CCU2D add_134_27 (.A0(\register[2][25] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][26] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24017), .COUT(n24018), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_27.INIT0 = 16'h5aaa;
    defparam add_134_27.INIT1 = 16'h5aaa;
    defparam add_134_27.INJECT1_0 = "NO";
    defparam add_134_27.INJECT1_1 = "NO";
    CCU2D add_134_25 (.A0(\register[2][23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24016), .COUT(n24017), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_25.INIT0 = 16'h5aaa;
    defparam add_134_25.INIT1 = 16'h5aaa;
    defparam add_134_25.INJECT1_0 = "NO";
    defparam add_134_25.INJECT1_1 = "NO";
    CCU2D add_134_23 (.A0(\register[2][21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24015), .COUT(n24016), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_23.INIT0 = 16'h5aaa;
    defparam add_134_23.INIT1 = 16'h5aaa;
    defparam add_134_23.INJECT1_0 = "NO";
    defparam add_134_23.INJECT1_1 = "NO";
    FD1P3IX read_size_i0_i1 (.D(n62), .SP(n12585), .CD(n26425), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n15_adj_243), .SP(n12585), .CD(n14798), 
            .CK(debug_c_c), .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n6739[0]), .SP(n12585), .CD(n8472), .CK(debug_c_c), 
            .Q(\read_value[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i0.GSR = "ENABLED";
    CCU2D add_134_21 (.A0(\register[2][19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24014), .COUT(n24015), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_21.INIT0 = 16'h5aaa;
    defparam add_134_21.INIT1 = 16'h5aaa;
    defparam add_134_21.INJECT1_0 = "NO";
    defparam add_134_21.INJECT1_1 = "NO";
    CCU2D add_134_19 (.A0(\register[2][17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24013), .COUT(n24014), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_19.INIT0 = 16'h5aaa;
    defparam add_134_19.INIT1 = 16'h5aaa;
    defparam add_134_19.INJECT1_0 = "NO";
    defparam add_134_19.INJECT1_1 = "NO";
    CCU2D add_134_17 (.A0(\register[2][15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24012), .COUT(n24013), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_17.INIT0 = 16'h5aaa;
    defparam add_134_17.INIT1 = 16'h5aaa;
    defparam add_134_17.INJECT1_0 = "NO";
    defparam add_134_17.INJECT1_1 = "NO";
    CCU2D add_134_15 (.A0(\register[2][13] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][14] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24011), .COUT(n24012), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_15.INIT0 = 16'h5aaa;
    defparam add_134_15.INIT1 = 16'h5aaa;
    defparam add_134_15.INJECT1_0 = "NO";
    defparam add_134_15.INJECT1_1 = "NO";
    CCU2D add_134_13 (.A0(\register[2][11] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][12] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24010), .COUT(n24011), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_13.INIT0 = 16'h5aaa;
    defparam add_134_13.INIT1 = 16'h5aaa;
    defparam add_134_13.INJECT1_0 = "NO";
    defparam add_134_13.INJECT1_1 = "NO";
    CCU2D add_134_11 (.A0(\register[2][9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][10] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24009), .COUT(n24010), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_11.INIT0 = 16'h5aaa;
    defparam add_134_11.INIT1 = 16'h5aaa;
    defparam add_134_11.INJECT1_0 = "NO";
    defparam add_134_11.INJECT1_1 = "NO";
    CCU2D add_134_9 (.A0(\register[2][7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][8] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24008), .COUT(n24009), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_9.INIT0 = 16'h5aaa;
    defparam add_134_9.INIT1 = 16'h5aaa;
    defparam add_134_9.INJECT1_0 = "NO";
    defparam add_134_9.INJECT1_1 = "NO";
    CCU2D add_134_7 (.A0(\register[2][5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24007), .COUT(n24008), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_7.INIT0 = 16'h5aaa;
    defparam add_134_7.INIT1 = 16'h5aaa;
    defparam add_134_7.INJECT1_0 = "NO";
    defparam add_134_7.INJECT1_1 = "NO";
    CCU2D add_134_5 (.A0(\register[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24006), .COUT(n24007), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_5.INIT0 = 16'h5aaa;
    defparam add_134_5.INIT1 = 16'h5aaa;
    defparam add_134_5.INJECT1_0 = "NO";
    defparam add_134_5.INJECT1_1 = "NO";
    CCU2D add_134_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24005), .COUT(n24006), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_3.INIT0 = 16'h5aaa;
    defparam add_134_3.INIT1 = 16'h5aaa;
    defparam add_134_3.INJECT1_0 = "NO";
    defparam add_134_3.INJECT1_1 = "NO";
    CCU2D add_134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24005), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_1.INIT0 = 16'hF000;
    defparam add_134_1.INIT1 = 16'h5555;
    defparam add_134_1.INJECT1_0 = "NO";
    defparam add_134_1.INJECT1_1 = "NO";
    LUT4 i13192_4_lut (.A(\register[2] [3]), .B(n15), .C(\register_addr[1] ), 
         .D(n4), .Z(n6739[3])) /* synthesis lut_function=(!(A (B ((D)+!C))+!A (B))) */ ;
    defparam i13192_4_lut.init = 16'h33b3;
    \ClockDividerP(factor=12000000)  uptime_div (.clk_1Hz(clk_1Hz), .debug_c_c(debug_c_c), 
            .n28477(n28477), .n2650(n2650), .GND_net(GND_net), .n26899(n26899)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(107[28] 109[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (clk_1Hz, debug_c_c, n28477, n2650, 
            GND_net, n26899) /* synthesis syn_module_defined=1 */ ;
    output clk_1Hz;
    input debug_c_c;
    input n28477;
    input n2650;
    input GND_net;
    output n26899;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7070;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n24296, n24295, n24294, n24293, n24292, n24291, n24290, 
        n24289, n24288, n24287, n24286, n24285, n24284, n24283, 
        n24282, n24281, n27, n24520, n25, n26, n24, n19, n32, 
        n28, n20, n29, n26_adj_466, n24224, n24223, n24222, n24221, 
        n24220, n24219, n24218, n24217, n24216, n24215, n24214, 
        n24213;
    
    FD1S3IX clk_o_14 (.D(n7070), .CK(debug_c_c), .CD(n28477), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2371__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2650), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i0.GSR = "ENABLED";
    CCU2D count_2371_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24296), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_33.INIT1 = 16'h0000;
    defparam count_2371_add_4_33.INJECT1_0 = "NO";
    defparam count_2371_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24295), .COUT(n24296), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_31.INJECT1_0 = "NO";
    defparam count_2371_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24294), .COUT(n24295), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_29.INJECT1_0 = "NO";
    defparam count_2371_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24293), .COUT(n24294), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_27.INJECT1_0 = "NO";
    defparam count_2371_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24292), .COUT(n24293), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_25.INJECT1_0 = "NO";
    defparam count_2371_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24291), .COUT(n24292), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_23.INJECT1_0 = "NO";
    defparam count_2371_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24290), .COUT(n24291), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_21.INJECT1_0 = "NO";
    defparam count_2371_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24289), .COUT(n24290), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_19.INJECT1_0 = "NO";
    defparam count_2371_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24288), .COUT(n24289), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_17.INJECT1_0 = "NO";
    defparam count_2371_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24287), .COUT(n24288), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_15.INJECT1_0 = "NO";
    defparam count_2371_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24286), .COUT(n24287), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_13.INJECT1_0 = "NO";
    defparam count_2371_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24285), .COUT(n24286), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_11.INJECT1_0 = "NO";
    defparam count_2371_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24284), .COUT(n24285), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_9.INJECT1_0 = "NO";
    defparam count_2371_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24283), .COUT(n24284), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_7.INJECT1_0 = "NO";
    defparam count_2371_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24282), .COUT(n24283), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_5.INJECT1_0 = "NO";
    defparam count_2371_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24281), .COUT(n24282), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2371_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2371_add_4_3.INJECT1_0 = "NO";
    defparam count_2371_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2371_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24281), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371_add_4_1.INIT0 = 16'hF000;
    defparam count_2371_add_4_1.INIT1 = 16'h0555;
    defparam count_2371_add_4_1.INJECT1_0 = "NO";
    defparam count_2371_add_4_1.INJECT1_1 = "NO";
    LUT4 i20300_4_lut (.A(n27), .B(n24520), .C(n25), .D(n26), .Z(n26899)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i20300_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n24520)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_466), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_396 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_396.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_397 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_397.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_466)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    FD1S3IX count_2371__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2650), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i1.GSR = "ENABLED";
    FD1S3IX count_2371__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2650), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i2.GSR = "ENABLED";
    FD1S3IX count_2371__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2650), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i3.GSR = "ENABLED";
    FD1S3IX count_2371__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2650), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i4.GSR = "ENABLED";
    FD1S3IX count_2371__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2650), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i5.GSR = "ENABLED";
    FD1S3IX count_2371__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2650), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i6.GSR = "ENABLED";
    FD1S3IX count_2371__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2650), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i7.GSR = "ENABLED";
    FD1S3IX count_2371__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2650), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i8.GSR = "ENABLED";
    FD1S3IX count_2371__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2650), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i9.GSR = "ENABLED";
    FD1S3IX count_2371__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i10.GSR = "ENABLED";
    FD1S3IX count_2371__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i11.GSR = "ENABLED";
    FD1S3IX count_2371__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i12.GSR = "ENABLED";
    FD1S3IX count_2371__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i13.GSR = "ENABLED";
    FD1S3IX count_2371__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i14.GSR = "ENABLED";
    FD1S3IX count_2371__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i15.GSR = "ENABLED";
    FD1S3IX count_2371__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i16.GSR = "ENABLED";
    FD1S3IX count_2371__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i17.GSR = "ENABLED";
    FD1S3IX count_2371__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i18.GSR = "ENABLED";
    FD1S3IX count_2371__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i19.GSR = "ENABLED";
    FD1S3IX count_2371__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i20.GSR = "ENABLED";
    FD1S3IX count_2371__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i21.GSR = "ENABLED";
    FD1S3IX count_2371__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i22.GSR = "ENABLED";
    FD1S3IX count_2371__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i23.GSR = "ENABLED";
    FD1S3IX count_2371__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i24.GSR = "ENABLED";
    FD1S3IX count_2371__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i25.GSR = "ENABLED";
    FD1S3IX count_2371__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i26.GSR = "ENABLED";
    FD1S3IX count_2371__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i27.GSR = "ENABLED";
    FD1S3IX count_2371__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i28.GSR = "ENABLED";
    FD1S3IX count_2371__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i29.GSR = "ENABLED";
    FD1S3IX count_2371__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i30.GSR = "ENABLED";
    FD1S3IX count_2371__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2650), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2371__i31.GSR = "ENABLED";
    CCU2D add_17801_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24224), 
          .S0(n7070));
    defparam add_17801_cout.INIT0 = 16'h0000;
    defparam add_17801_cout.INIT1 = 16'h0000;
    defparam add_17801_cout.INJECT1_0 = "NO";
    defparam add_17801_cout.INJECT1_1 = "NO";
    CCU2D add_17801_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24223), .COUT(n24224));
    defparam add_17801_24.INIT0 = 16'h5555;
    defparam add_17801_24.INIT1 = 16'h5555;
    defparam add_17801_24.INJECT1_0 = "NO";
    defparam add_17801_24.INJECT1_1 = "NO";
    CCU2D add_17801_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24222), .COUT(n24223));
    defparam add_17801_22.INIT0 = 16'h5555;
    defparam add_17801_22.INIT1 = 16'h5555;
    defparam add_17801_22.INJECT1_0 = "NO";
    defparam add_17801_22.INJECT1_1 = "NO";
    CCU2D add_17801_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24221), .COUT(n24222));
    defparam add_17801_20.INIT0 = 16'h5555;
    defparam add_17801_20.INIT1 = 16'h5555;
    defparam add_17801_20.INJECT1_0 = "NO";
    defparam add_17801_20.INJECT1_1 = "NO";
    CCU2D add_17801_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24220), .COUT(n24221));
    defparam add_17801_18.INIT0 = 16'h5555;
    defparam add_17801_18.INIT1 = 16'h5555;
    defparam add_17801_18.INJECT1_0 = "NO";
    defparam add_17801_18.INJECT1_1 = "NO";
    CCU2D add_17801_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24219), .COUT(n24220));
    defparam add_17801_16.INIT0 = 16'h5aaa;
    defparam add_17801_16.INIT1 = 16'h5555;
    defparam add_17801_16.INJECT1_0 = "NO";
    defparam add_17801_16.INJECT1_1 = "NO";
    CCU2D add_17801_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24218), .COUT(n24219));
    defparam add_17801_14.INIT0 = 16'h5aaa;
    defparam add_17801_14.INIT1 = 16'h5555;
    defparam add_17801_14.INJECT1_0 = "NO";
    defparam add_17801_14.INJECT1_1 = "NO";
    CCU2D add_17801_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24217), .COUT(n24218));
    defparam add_17801_12.INIT0 = 16'h5555;
    defparam add_17801_12.INIT1 = 16'h5aaa;
    defparam add_17801_12.INJECT1_0 = "NO";
    defparam add_17801_12.INJECT1_1 = "NO";
    CCU2D add_17801_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24216), .COUT(n24217));
    defparam add_17801_10.INIT0 = 16'h5aaa;
    defparam add_17801_10.INIT1 = 16'h5aaa;
    defparam add_17801_10.INJECT1_0 = "NO";
    defparam add_17801_10.INJECT1_1 = "NO";
    CCU2D add_17801_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24215), .COUT(n24216));
    defparam add_17801_8.INIT0 = 16'h5555;
    defparam add_17801_8.INIT1 = 16'h5aaa;
    defparam add_17801_8.INJECT1_0 = "NO";
    defparam add_17801_8.INJECT1_1 = "NO";
    CCU2D add_17801_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24214), .COUT(n24215));
    defparam add_17801_6.INIT0 = 16'h5555;
    defparam add_17801_6.INIT1 = 16'h5555;
    defparam add_17801_6.INJECT1_0 = "NO";
    defparam add_17801_6.INJECT1_1 = "NO";
    CCU2D add_17801_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24213), .COUT(n24214));
    defparam add_17801_4.INIT0 = 16'h5aaa;
    defparam add_17801_4.INIT1 = 16'h5aaa;
    defparam add_17801_4.INJECT1_0 = "NO";
    defparam add_17801_4.INJECT1_1 = "NO";
    CCU2D add_17801_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24213));
    defparam add_17801_2.INIT0 = 16'h7000;
    defparam add_17801_2.INIT1 = 16'h5555;
    defparam add_17801_2.INJECT1_0 = "NO";
    defparam add_17801_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module SabertoothSerialPeripheral
//

module SabertoothSerialPeripheral (\register[1] , debug_c_c, n282, n28477, 
            \databus[6] , \databus[5] , \databus[4] , \databus[3] , 
            \databus[2] , \register[1][1] , \databus[1] , \databus[0] , 
            \register[0] , \register[0][4] , \register[0][1] , \read_size[0] , 
            n28425, \select[2] , read_value, rw, n64, n28415, \register_addr[0] , 
            n28560, n4, n28537, n19865, n22, \reset_count[14] , 
            n82, \register_addr[2] , n28440, n28443, \state[0] , GND_net, 
            n12, \state[1] , n28405, n6599, n17488, n21, n7, n19338, 
            n25733, n28505, n962, n17481, n89, n41, n32, n87, 
            n31, n86, n30, n88, n29, n28, n5069, n5068, n5067, 
            n5066, n5065, n28504, n28506, state, n27784, n13009, 
            n24633, n19370, \reset_count[11] , \reset_count[8] , n24551, 
            n26512, \reset_count[7] , n26556, motor_pwm_l_c, n27404, 
            n46, n7_adj_237, \reset_count[6] , \reset_count[5] , \reset_count[4] , 
            n47, n2736, select_clk, n16717, n7591, n28406, n26896) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\register[1] ;
    input debug_c_c;
    input n282;
    input n28477;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    output \register[1][1] ;
    input \databus[1] ;
    input \databus[0] ;
    output [7:0]\register[0] ;
    output \register[0][4] ;
    output \register[0][1] ;
    output \read_size[0] ;
    input n28425;
    input \select[2] ;
    output [7:0]read_value;
    input rw;
    output n64;
    input n28415;
    input \register_addr[0] ;
    output n28560;
    output n4;
    input n28537;
    output n19865;
    output n22;
    input \reset_count[14] ;
    input n82;
    input \register_addr[2] ;
    input n28440;
    output n28443;
    output \state[0] ;
    input GND_net;
    input n12;
    output \state[1] ;
    input n28405;
    input n6599;
    output n17488;
    input n21;
    output n7;
    input n19338;
    input n25733;
    input n28505;
    output n962;
    input n17481;
    output n89;
    output n41;
    output n32;
    output n87;
    output n31;
    output n86;
    output n30;
    output n88;
    output n29;
    output n28;
    input n5069;
    input n5068;
    input n5067;
    input n5066;
    input n5065;
    input n28504;
    input n28506;
    output [3:0]state;
    input n27784;
    input n13009;
    input n24633;
    input n19370;
    input \reset_count[11] ;
    input \reset_count[8] ;
    input n24551;
    output n26512;
    input \reset_count[7] ;
    output n26556;
    output motor_pwm_l_c;
    input n27404;
    output n46;
    input n7_adj_237;
    input \reset_count[6] ;
    input \reset_count[5] ;
    input \reset_count[4] ;
    output n47;
    input n2736;
    output select_clk;
    input n16717;
    output n7591;
    output n28406;
    output n26896;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n12620;
    wire [7:0]\register[1]_c ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n28408, n19955;
    wire [7:0]\register[0]_c ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n28407, n2606, prev_select, n8476;
    wire [7:0]n5133;
    
    wire n28575, n28561, n28472, n28503, n17519, n28562, n28507, 
        n28473, n17494, n19561, n24509, n28446;
    
    FD1P3AX register_0__i16 (.D(n282), .SP(n12620), .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n28408), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[1]_c [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n28408), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[1]_c [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n28408), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[1]_c [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n28408), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[1]_c [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n28408), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[1]_c [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n28408), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[1][1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n28408), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[1]_c [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n282), .SP(n19955), .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n28407), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[0]_c [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n28407), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[0]_c [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n28407), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[0][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n28407), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[0]_c [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n28407), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[0]_c [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n28407), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[0][1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i2.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n28425), .SP(n2606), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n28407), .PD(n28477), 
            .CK(debug_c_c), .Q(\register[0]_c [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam prev_select_138.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n5133[0]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n5133[7]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n5133[6]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n5133[5]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5133[4]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5133[3]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n5133[2]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n5133[1]), .SP(n2606), .CD(n8476), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i16_2_lut (.A(\select[2] ), .B(rw), .Z(n64)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam i16_2_lut.init = 16'h8888;
    LUT4 i20319_2_lut_3_lut_4_lut (.A(n28575), .B(n28415), .C(n28477), 
         .D(\register_addr[0] ), .Z(n19955)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam i20319_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n28575), .B(n28415), .C(n28477), .D(\register_addr[0] ), 
         .Z(n12620)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 i1_2_lut_rep_439 (.A(\register[0]_c [3]), .B(\register[0]_c [2]), 
         .Z(n28560)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_2_lut_rep_439.init = 16'h8888;
    LUT4 i1_2_lut_rep_351_3_lut_4_lut (.A(\register[0]_c [3]), .B(\register[0]_c [2]), 
         .C(n28561), .D(\register[0][1] ), .Z(n28472)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_2_lut_rep_351_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_382_3_lut (.A(\register[0]_c [3]), .B(\register[0]_c [2]), 
         .C(\register[0][1] ), .Z(n28503)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_2_lut_rep_382_3_lut.init = 16'h8080;
    LUT4 i13_2_lut_3_lut_4_lut (.A(\register[0]_c [3]), .B(\register[0]_c [2]), 
         .C(\register[0][4] ), .D(\register[0][1] ), .Z(n17519)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i13_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_rep_440 (.A(\register[0]_c [6]), .B(\register[0]_c [5]), 
         .Z(n28561)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_2_lut_rep_440.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(\register[0]_c [6]), .B(\register[0]_c [5]), 
         .C(\register[0]_c [0]), .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_441 (.A(\register[1]_c [2]), .B(\register[1][1] ), 
         .Z(n28562)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_2_lut_rep_441.init = 16'h8888;
    LUT4 i1_2_lut_rep_386_3_lut (.A(\register[1]_c [2]), .B(\register[1][1] ), 
         .C(\register[1]_c [3]), .Z(n28507)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_2_lut_rep_386_3_lut.init = 16'h8080;
    LUT4 i5523_2_lut_rep_352_3_lut_4_lut (.A(\register[1]_c [2]), .B(\register[1][1] ), 
         .C(\register[1]_c [4]), .D(\register[1]_c [3]), .Z(n28473)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i5523_2_lut_rep_352_3_lut_4_lut.init = 16'h8000;
    LUT4 i11499_3_lut_4_lut (.A(\register[0][1] ), .B(n28560), .C(\register[0][4] ), 
         .D(\register[0]_c [5]), .Z(n17494)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i11499_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_4_lut_4_lut (.A(\register[1][1] ), .B(n28537), .C(n19865), 
         .D(\register[1]_c [2]), .Z(n22)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i1_4_lut_4_lut.init = 16'hf1e2;
    LUT4 i1_4_lut_4_lut_adj_395 (.A(\register[1] [7]), .B(n28537), .C(n19561), 
         .D(n24509), .Z(n19865)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i1_4_lut_4_lut_adj_395.init = 16'h2000;
    LUT4 i5527_2_lut_rep_325_3_lut_4_lut (.A(\register[1]_c [3]), .B(n28562), 
         .C(\register[1]_c [5]), .D(\register[1]_c [4]), .Z(n28446)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i5527_2_lut_rep_325_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_454 (.A(\select[2] ), .B(prev_select), .Z(n28575)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_rep_454.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\select[2] ), .B(prev_select), .C(\reset_count[14] ), 
         .D(n82), .Z(n2606)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i3_4_lut (.A(\register[1]_c [3]), .B(\register[1]_c [2]), .C(\register[1]_c [5]), 
         .D(\register[1]_c [6]), .Z(n24509)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2_4_lut (.A(n28575), .B(n28477), .C(\register_addr[2] ), .D(n28440), 
         .Z(n8476)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i2_4_lut.init = 16'h2220;
    LUT4 mux_1721_Mux_0_i1_3_lut (.A(\register[0]_c [0]), .B(\register[1]_c [0]), 
         .C(\register_addr[0] ), .Z(n5133[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1721_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1721_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n5133[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1721_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1721_Mux_6_i1_3_lut (.A(\register[0]_c [6]), .B(\register[1]_c [6]), 
         .C(\register_addr[0] ), .Z(n5133[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1721_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1721_Mux_4_i1_3_lut (.A(\register[0][4] ), .B(\register[1]_c [4]), 
         .C(\register_addr[0] ), .Z(n5133[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1721_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 i11694_3_lut (.A(\register[0]_c [3]), .B(\register[1]_c [3]), .C(\register_addr[0] ), 
         .Z(n5133[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11694_3_lut.init = 16'hcaca;
    LUT4 i11695_3_lut (.A(\register[0]_c [2]), .B(\register[1]_c [2]), .C(\register_addr[0] ), 
         .Z(n5133[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11695_3_lut.init = 16'hcaca;
    LUT4 i11698_3_lut (.A(\register[0][1] ), .B(\register[1][1] ), .C(\register_addr[0] ), 
         .Z(n5133[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11698_3_lut.init = 16'hcaca;
    LUT4 i20322_2_lut_rep_286_3_lut_4_lut (.A(rw), .B(n28425), .C(\register_addr[0] ), 
         .D(n28575), .Z(n28407)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i20322_2_lut_rep_286_3_lut_4_lut.init = 16'h0400;
    LUT4 i4262_2_lut_rep_287_3_lut_4_lut (.A(rw), .B(n28425), .C(\register_addr[0] ), 
         .D(n28575), .Z(n28408)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i4262_2_lut_rep_287_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_3_lut_rep_322_4_lut (.A(n28503), .B(n28561), .C(\register[0][4] ), 
         .D(n28537), .Z(n28443)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i1_3_lut_rep_322_4_lut.init = 16'hff80;
    SabertoothSerial sserial (.\state[0] (\state[0] ), .debug_c_c(debug_c_c), 
            .GND_net(GND_net), .n12(n12), .\state[1] (\state[1] ), .n28405(n28405), 
            .n6599(n6599), .n28443(n28443), .n17488(n17488), .n21(n21), 
            .n7(n7), .n19338(n19338), .n25733(n25733), .n28505(n28505), 
            .\register[1][7] (\register[1] [7]), .n28537(n28537), .n962(n962), 
            .n17481(n17481), .\register[0] ({\register[0] [7], \register[0]_c [6:5], 
            \register[0][4] , \register[0]_c [3:2], \register[0][1] , 
            \register[0]_c [0]}), .n28472(n28472), .\register[1][0] (\register[1]_c [0]), 
            .\register[1][4] (\register[1]_c [4]), .n19561(n19561), .n28562(n28562), 
            .\register[1][3] (\register[1]_c [3]), .n89(n89), .n41(n41), 
            .n32(n32), .\register[1][5] (\register[1]_c [5]), .n28473(n28473), 
            .n87(n87), .n17494(n17494), .n31(n31), .\register[1][6] (\register[1]_c [6]), 
            .n28446(n28446), .n86(n86), .n30(n30), .n28560(n28560), 
            .n28507(n28507), .n88(n88), .n17519(n17519), .n29(n29), 
            .n28(n28), .n5069(n5069), .\register_addr[0] (\register_addr[0] ), 
            .n5136(n5133[5]), .n5068(n5068), .n5067(n5067), .n5066(n5066), 
            .n5065(n5065), .n28504(n28504), .n19865(n19865), .n28506(n28506), 
            .n28477(n28477), .state({state}), .n27784(n27784), .n13009(n13009), 
            .n24633(n24633), .n19370(n19370), .\reset_count[11] (\reset_count[11] ), 
            .\reset_count[8] (\reset_count[8] ), .n24551(n24551), .n26512(n26512), 
            .\reset_count[7] (\reset_count[7] ), .n26556(n26556), .motor_pwm_l_c(motor_pwm_l_c), 
            .n27404(n27404), .n46(n46), .n7_adj_234(n7_adj_237), .\reset_count[14] (\reset_count[14] ), 
            .n82(n82), .\reset_count[6] (\reset_count[6] ), .\reset_count[5] (\reset_count[5] ), 
            .\reset_count[4] (\reset_count[4] ), .n47(n47), .n2736(n2736), 
            .select_clk(select_clk), .n16717(n16717), .n7591(n7591), .n28406(n28406), 
            .n26896(n26896)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(142[19] 147[34])
    
endmodule
//
// Verilog Description of module SabertoothSerial
//

module SabertoothSerial (\state[0] , debug_c_c, GND_net, n12, \state[1] , 
            n28405, n6599, n28443, n17488, n21, n7, n19338, n25733, 
            n28505, \register[1][7] , n28537, n962, n17481, \register[0] , 
            n28472, \register[1][0] , \register[1][4] , n19561, n28562, 
            \register[1][3] , n89, n41, n32, \register[1][5] , n28473, 
            n87, n17494, n31, \register[1][6] , n28446, n86, n30, 
            n28560, n28507, n88, n17519, n29, n28, n5069, \register_addr[0] , 
            n5136, n5068, n5067, n5066, n5065, n28504, n19865, 
            n28506, n28477, state, n27784, n13009, n24633, n19370, 
            \reset_count[11] , \reset_count[8] , n24551, n26512, \reset_count[7] , 
            n26556, motor_pwm_l_c, n27404, n46, n7_adj_234, \reset_count[14] , 
            n82, \reset_count[6] , \reset_count[5] , \reset_count[4] , 
            n47, n2736, select_clk, n16717, n7591, n28406, n26896) /* synthesis syn_module_defined=1 */ ;
    output \state[0] ;
    input debug_c_c;
    input GND_net;
    input n12;
    output \state[1] ;
    input n28405;
    input n6599;
    input n28443;
    output n17488;
    input n21;
    output n7;
    input n19338;
    input n25733;
    input n28505;
    input \register[1][7] ;
    input n28537;
    output n962;
    input n17481;
    input [7:0]\register[0] ;
    input n28472;
    input \register[1][0] ;
    input \register[1][4] ;
    output n19561;
    input n28562;
    input \register[1][3] ;
    output n89;
    output n41;
    output n32;
    input \register[1][5] ;
    input n28473;
    output n87;
    input n17494;
    output n31;
    input \register[1][6] ;
    input n28446;
    output n86;
    output n30;
    input n28560;
    input n28507;
    output n88;
    input n17519;
    output n29;
    output n28;
    input n5069;
    input \register_addr[0] ;
    output n5136;
    input n5068;
    input n5067;
    input n5066;
    input n5065;
    input n28504;
    input n19865;
    input n28506;
    input n28477;
    output [3:0]state;
    input n27784;
    input n13009;
    input n24633;
    input n19370;
    input \reset_count[11] ;
    input \reset_count[8] ;
    input n24551;
    output n26512;
    input \reset_count[7] ;
    output n26556;
    output motor_pwm_l_c;
    input n27404;
    output n46;
    input n7_adj_234;
    input \reset_count[14] ;
    input n82;
    input \reset_count[6] ;
    input \reset_count[5] ;
    input \reset_count[4] ;
    output n47;
    input n2736;
    output select_clk;
    input n16717;
    output n7591;
    output n28406;
    output n26896;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(16[12:19])
    
    wire n28404;
    wire [7:0]n5062;
    
    wire n27723, n27725;
    wire [31:0]n59;
    
    wire n9285, n27726, n9034, n17524, n17515, n4, n17528, n27727;
    
    FD1S3IX state__i0 (.D(n12), .CK(debug_c_c), .CD(GND_net), .Q(\state[0] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n5062[0]), .SP(n28404), .CK(debug_c_c), 
            .Q(tx_data[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1P3IX state__i1 (.D(n6599), .SP(n28405), .CD(GND_net), .CK(debug_c_c), 
            .Q(\state[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 n27724_bdd_2_lut_3_lut (.A(n27723), .B(n28443), .C(n17488), .Z(n27725)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam n27724_bdd_2_lut_3_lut.init = 16'h0808;
    PFUMX mux_1714_i7 (.BLUT(n59[6]), .ALUT(n21), .C0(n7), .Z(n5062[6]));
    PFUMX mux_1714_i1 (.BLUT(n19338), .ALUT(n25733), .C0(n7), .Z(n5062[0]));
    LUT4 n17488_bdd_4_lut_20631 (.A(n9285), .B(n28505), .C(\register[1][7] ), 
         .D(n28537), .Z(n27726)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam n17488_bdd_4_lut_20631.init = 16'hffdf;
    FD1P3AX send_27 (.D(n9034), .SP(n28405), .CK(debug_c_c), .Q(n962));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam send_27.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\state[0] ), .B(\state[1] ), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut (.A(n17481), .B(n28537), .C(\register[0] [0]), .D(n28472), 
         .Z(n17488)) /* synthesis lut_function=(A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(494[7:19])
    defparam i1_4_lut.init = 16'ha888;
    LUT4 i13350_2_lut (.A(\register[1][0] ), .B(\register[1][4] ), .Z(n19561)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13350_2_lut.init = 16'h8888;
    LUT4 i13640_4_lut (.A(n28562), .B(n28505), .C(n28537), .D(\register[1][3] ), 
         .Z(n89)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i13640_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_389 (.A(n28537), .B(n41), .C(n17488), .D(n17524), 
         .Z(n32)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_389.init = 16'h3130;
    LUT4 n9235_bdd_4_lut_20692 (.A(\register[0] [7]), .B(\state[1] ), .C(\state[0] ), 
         .D(n28537), .Z(n27723)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam n9235_bdd_4_lut_20692.init = 16'h0002;
    LUT4 i11529_3_lut (.A(\register[0] [3]), .B(\register[0] [1]), .C(\register[0] [2]), 
         .Z(n17524)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    defparam i11529_3_lut.init = 16'h6a6a;
    LUT4 i41_2_lut (.A(\state[0] ), .B(\state[1] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i41_2_lut.init = 16'heeee;
    LUT4 i13642_4_lut (.A(\register[1][5] ), .B(n28505), .C(n28537), .D(n28473), 
         .Z(n87)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i13642_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_390 (.A(n28537), .B(n41), .C(n17488), .D(n17494), 
         .Z(n31)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_390.init = 16'h3130;
    LUT4 i13643_4_lut (.A(\register[1][6] ), .B(n28505), .C(n28537), .D(n28446), 
         .Z(n86)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i13643_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_391 (.A(n28537), .B(n41), .C(n17488), .D(n17515), 
         .Z(n30)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_391.init = 16'h3130;
    LUT4 i13181_4_lut (.A(\register[0] [6]), .B(\register[0] [1]), .C(n28560), 
         .D(n4), .Z(n17515)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam i13181_4_lut.init = 16'h6aaa;
    LUT4 i1_2_lut_adj_392 (.A(\register[0] [4]), .B(\register[0] [5]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    defparam i1_2_lut_adj_392.init = 16'h8888;
    LUT4 i13641_4_lut (.A(\register[1][4] ), .B(n28505), .C(n28537), .D(n28507), 
         .Z(n88)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i13641_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_393 (.A(n28537), .B(n41), .C(n17488), .D(n17519), 
         .Z(n29)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_393.init = 16'h3130;
    LUT4 i1_4_lut_adj_394 (.A(n28537), .B(n41), .C(n17488), .D(n17528), 
         .Z(n28)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_394.init = 16'h3130;
    LUT4 i15_2_lut (.A(\register[0] [1]), .B(\register[0] [2]), .Z(n17528)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    defparam i15_2_lut.init = 16'h6666;
    FD1P3AX tx_data_i0_i1 (.D(n5069), .SP(n28404), .CK(debug_c_c), .Q(tx_data[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    PFUMX i20629 (.BLUT(n27726), .ALUT(n27725), .C0(n7), .Z(n27727));
    LUT4 i11559_3_lut (.A(\register[0] [5]), .B(\register[1][5] ), .C(\register_addr[0] ), 
         .Z(n5136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11559_3_lut.init = 16'hcaca;
    FD1P3AX tx_data_i0_i2 (.D(n5068), .SP(n28404), .CK(debug_c_c), .Q(tx_data[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n5067), .SP(n28404), .CK(debug_c_c), .Q(tx_data[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n5066), .SP(n28404), .CK(debug_c_c), .Q(tx_data[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i5 (.D(n5065), .SP(n28404), .CK(debug_c_c), .Q(tx_data[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i6 (.D(n5062[6]), .SP(n28404), .CK(debug_c_c), 
            .Q(tx_data[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i7 (.D(n27727), .SP(n28404), .CK(debug_c_c), .Q(tx_data[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i13644_3_lut_4_lut (.A(n28504), .B(n19865), .C(n9285), .D(n28506), 
         .Z(n59[6])) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;
    defparam i13644_3_lut_4_lut.init = 16'h8ff8;
    LUT4 i10742_1_lut (.A(\state[0] ), .Z(n9034)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i10742_1_lut.init = 16'h5555;
    LUT4 i13750_3_lut_4_lut (.A(\register[1][5] ), .B(n28473), .C(n28537), 
         .D(\register[1][6] ), .Z(n9285)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i13750_3_lut_4_lut.init = 16'hf8f0;
    \UARTTransmitter(baud_div=1250)  sender (.n28477(n28477), .state({state}), 
            .n27784(n27784), .n13009(n13009), .n24633(n24633), .n19370(n19370), 
            .\reset_count[11] (\reset_count[11] ), .\reset_count[8] (\reset_count[8] ), 
            .n24551(n24551), .n26512(n26512), .tx_data({tx_data}), .\reset_count[7] (\reset_count[7] ), 
            .n26556(n26556), .motor_pwm_l_c(motor_pwm_l_c), .n27404(n27404), 
            .n46(n46), .n7(n7_adj_234), .n962(n962), .\reset_count[14] (\reset_count[14] ), 
            .n82(n82), .\reset_count[6] (\reset_count[6] ), .\reset_count[5] (\reset_count[5] ), 
            .\reset_count[4] (\reset_count[4] ), .n47(n47), .GND_net(GND_net), 
            .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(63[26] 67[47])
    \ClockDividerP(factor=12000)  baud_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .n2736(n2736), .select_clk(select_clk), .n16717(n16717), .n7591(n7591), 
            .n28406(n28406), .\state[0] (\state[0] ), .n28477(n28477), 
            .n28404(n28404), .n26896(n26896)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(21[25] 23[48])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=1250) 
//

module \UARTTransmitter(baud_div=1250)  (n28477, state, n27784, n13009, 
            n24633, n19370, \reset_count[11] , \reset_count[8] , n24551, 
            n26512, tx_data, \reset_count[7] , n26556, motor_pwm_l_c, 
            n27404, n46, n7, n962, \reset_count[14] , n82, \reset_count[6] , 
            \reset_count[5] , \reset_count[4] , n47, GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input n28477;
    output [3:0]state;
    input n27784;
    input n13009;
    input n24633;
    input n19370;
    input \reset_count[11] ;
    input \reset_count[8] ;
    input n24551;
    output n26512;
    input [7:0]tx_data;
    input \reset_count[7] ;
    output n26556;
    output motor_pwm_l_c;
    input n27404;
    output n46;
    input n7;
    input n962;
    input \reset_count[14] ;
    input n82;
    input \reset_count[6] ;
    input \reset_count[5] ;
    input \reset_count[4] ;
    output n47;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n26770, n26340, n7_c, n10, n104, n26856, n26857, n26858;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n8397, n2, n26341;
    
    LUT4 i1_4_lut (.A(n28477), .B(state[1]), .C(n26770), .D(state[0]), 
         .Z(n26340)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0104;
    FD1S3IX state__i0 (.D(n27784), .CK(bclk), .CD(n28477), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 i20076_2_lut (.A(state[2]), .B(state[3]), .Z(n26770)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20076_2_lut.init = 16'h8888;
    FD1P3AX state__i3 (.D(n24633), .SP(n13009), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_386 (.A(n19370), .B(\reset_count[11] ), .C(\reset_count[8] ), 
         .D(n24551), .Z(n26512)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_386.init = 16'h8880;
    PFUMX Mux_22_i15 (.BLUT(n7_c), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;
    PFUMX i20162 (.BLUT(n26856), .ALUT(n26857), .C0(state[1]), .Z(n26858));
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n8397), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\reset_count[8] ), .B(\reset_count[7] ), .Z(n26556)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3JX tx_35 (.D(n104), .SP(n27404), .PD(n28477), .CK(bclk), .Q(motor_pwm_l_c)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n26858), .C(state[2]), .D(state[1]), 
         .Z(n7_c)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i13694_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i13694_4_lut.init = 16'hfcee;
    LUT4 i20160_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n26856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20160_3_lut.init = 16'hcaca;
    LUT4 i20161_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n26857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20161_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_387 (.A(state[1]), .B(state[0]), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_2_lut_adj_387.init = 16'h8888;
    FD1P3AX state__i1 (.D(n26340), .SP(n13009), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX state__i2 (.D(n7), .SP(n13009), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n8397), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n8397), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n8397), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n8397), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n8397), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n8397), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n8397), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(state[3]), .B(n962), .C(\reset_count[14] ), .D(n26341), 
         .Z(n8397)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut.init = 16'h4000;
    LUT4 i3_4_lut_adj_388 (.A(n82), .B(state[0]), .C(state[2]), .D(state[1]), 
         .Z(n26341)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_388.init = 16'h0002;
    LUT4 i1_3_lut (.A(\reset_count[6] ), .B(\reset_count[5] ), .C(\reset_count[4] ), 
         .Z(n47)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i1_3_lut.init = 16'ha8a8;
    \ClockDividerP(factor=1250)  baud_gen (.GND_net(GND_net), .bclk(bclk), 
            .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=1250) 
//

module \ClockDividerP(factor=1250)  (GND_net, bclk, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output bclk;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24392;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n102;
    
    wire n24391, n24390, n24389, n24388, n24387, n24386, n24385, 
        n24384, n24383, n24382, n24381, n24380, n24379, n24378, 
        n24377, n26961, n45, n52, n46, n14872, n50, n42, n48, 
        n38, n44, n30, n26774, n7626, n24476, n24475, n24474, 
        n24473, n24472, n24471, n24470, n24469, n24468, n24467, 
        n24466, n24465, n24464, n24463, n24462;
    
    CCU2D count_2379_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24392), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_33.INIT1 = 16'h0000;
    defparam count_2379_add_4_33.INJECT1_0 = "NO";
    defparam count_2379_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24391), .COUT(n24392), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_31.INJECT1_0 = "NO";
    defparam count_2379_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24390), .COUT(n24391), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_29.INJECT1_0 = "NO";
    defparam count_2379_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24389), .COUT(n24390), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_27.INJECT1_0 = "NO";
    defparam count_2379_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24388), .COUT(n24389), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_25.INJECT1_0 = "NO";
    defparam count_2379_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24387), .COUT(n24388), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_23.INJECT1_0 = "NO";
    defparam count_2379_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24386), .COUT(n24387), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_21.INJECT1_0 = "NO";
    defparam count_2379_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24385), .COUT(n24386), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_19.INJECT1_0 = "NO";
    defparam count_2379_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24384), .COUT(n24385), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_17.INJECT1_0 = "NO";
    defparam count_2379_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24383), .COUT(n24384), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_15.INJECT1_0 = "NO";
    defparam count_2379_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24382), .COUT(n24383), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_13.INJECT1_0 = "NO";
    defparam count_2379_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24381), .COUT(n24382), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_11.INJECT1_0 = "NO";
    defparam count_2379_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24380), .COUT(n24381), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_9.INJECT1_0 = "NO";
    defparam count_2379_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24379), .COUT(n24380), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_7.INJECT1_0 = "NO";
    defparam count_2379_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24378), .COUT(n24379), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_5.INJECT1_0 = "NO";
    defparam count_2379_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24377), .COUT(n24378), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2379_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2379_add_4_3.INJECT1_0 = "NO";
    defparam count_2379_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2379_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24377), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379_add_4_1.INIT0 = 16'hF000;
    defparam count_2379_add_4_1.INIT1 = 16'h0555;
    defparam count_2379_add_4_1.INJECT1_0 = "NO";
    defparam count_2379_add_4_1.INJECT1_1 = "NO";
    LUT4 i20364_4_lut (.A(n26961), .B(n45), .C(n52), .D(n46), .Z(n14872)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20364_4_lut.init = 16'h0002;
    LUT4 i20362_4_lut (.A(count[13]), .B(n50), .C(n42), .D(count[3]), 
         .Z(n26961)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20362_4_lut.init = 16'h0001;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n45)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(count[30]), .B(n48), .C(n38), .D(count[14]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(count[24]), .B(count[4]), .C(count[1]), .D(count[27]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(count[28]), .B(n44), .C(n30), .D(count[18]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(count[31]), .B(count[5]), .C(n26774), .D(count[6]), 
         .Z(n42)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i14_4_lut.init = 16'hbfff;
    LUT4 i16_4_lut (.A(count[16]), .B(count[21]), .C(count[11]), .D(count[25]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[2]), .B(count[8]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(count[20]), .B(count[23]), .C(count[15]), .D(count[29]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(count[19]), .B(count[22]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i20080_3_lut (.A(count[10]), .B(count[0]), .C(count[7]), .Z(n26774)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i20080_3_lut.init = 16'h8080;
    FD1S3AX clk_o_14 (.D(n7626), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2379__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i0.GSR = "ENABLED";
    CCU2D add_17802_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24476), 
          .S1(n7626));
    defparam add_17802_32.INIT0 = 16'h5555;
    defparam add_17802_32.INIT1 = 16'h0000;
    defparam add_17802_32.INJECT1_0 = "NO";
    defparam add_17802_32.INJECT1_1 = "NO";
    CCU2D add_17802_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24475), .COUT(n24476));
    defparam add_17802_30.INIT0 = 16'h5555;
    defparam add_17802_30.INIT1 = 16'h5555;
    defparam add_17802_30.INJECT1_0 = "NO";
    defparam add_17802_30.INJECT1_1 = "NO";
    CCU2D add_17802_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24474), .COUT(n24475));
    defparam add_17802_28.INIT0 = 16'h5555;
    defparam add_17802_28.INIT1 = 16'h5555;
    defparam add_17802_28.INJECT1_0 = "NO";
    defparam add_17802_28.INJECT1_1 = "NO";
    CCU2D add_17802_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24473), .COUT(n24474));
    defparam add_17802_26.INIT0 = 16'h5555;
    defparam add_17802_26.INIT1 = 16'h5555;
    defparam add_17802_26.INJECT1_0 = "NO";
    defparam add_17802_26.INJECT1_1 = "NO";
    CCU2D add_17802_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24472), .COUT(n24473));
    defparam add_17802_24.INIT0 = 16'h5555;
    defparam add_17802_24.INIT1 = 16'h5555;
    defparam add_17802_24.INJECT1_0 = "NO";
    defparam add_17802_24.INJECT1_1 = "NO";
    CCU2D add_17802_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24471), .COUT(n24472));
    defparam add_17802_22.INIT0 = 16'h5555;
    defparam add_17802_22.INIT1 = 16'h5555;
    defparam add_17802_22.INJECT1_0 = "NO";
    defparam add_17802_22.INJECT1_1 = "NO";
    CCU2D add_17802_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24470), .COUT(n24471));
    defparam add_17802_20.INIT0 = 16'h5555;
    defparam add_17802_20.INIT1 = 16'h5555;
    defparam add_17802_20.INJECT1_0 = "NO";
    defparam add_17802_20.INJECT1_1 = "NO";
    CCU2D add_17802_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24469), .COUT(n24470));
    defparam add_17802_18.INIT0 = 16'h5555;
    defparam add_17802_18.INIT1 = 16'h5555;
    defparam add_17802_18.INJECT1_0 = "NO";
    defparam add_17802_18.INJECT1_1 = "NO";
    CCU2D add_17802_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24468), .COUT(n24469));
    defparam add_17802_16.INIT0 = 16'h5555;
    defparam add_17802_16.INIT1 = 16'h5555;
    defparam add_17802_16.INJECT1_0 = "NO";
    defparam add_17802_16.INJECT1_1 = "NO";
    CCU2D add_17802_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24467), .COUT(n24468));
    defparam add_17802_14.INIT0 = 16'h5555;
    defparam add_17802_14.INIT1 = 16'h5555;
    defparam add_17802_14.INJECT1_0 = "NO";
    defparam add_17802_14.INJECT1_1 = "NO";
    CCU2D add_17802_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24466), .COUT(n24467));
    defparam add_17802_12.INIT0 = 16'h5555;
    defparam add_17802_12.INIT1 = 16'h5555;
    defparam add_17802_12.INJECT1_0 = "NO";
    defparam add_17802_12.INJECT1_1 = "NO";
    CCU2D add_17802_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24465), .COUT(n24466));
    defparam add_17802_10.INIT0 = 16'h5aaa;
    defparam add_17802_10.INIT1 = 16'h5555;
    defparam add_17802_10.INJECT1_0 = "NO";
    defparam add_17802_10.INJECT1_1 = "NO";
    CCU2D add_17802_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24464), 
          .COUT(n24465));
    defparam add_17802_8.INIT0 = 16'h5555;
    defparam add_17802_8.INIT1 = 16'h5555;
    defparam add_17802_8.INJECT1_0 = "NO";
    defparam add_17802_8.INJECT1_1 = "NO";
    CCU2D add_17802_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24463), 
          .COUT(n24464));
    defparam add_17802_6.INIT0 = 16'h5aaa;
    defparam add_17802_6.INIT1 = 16'h5aaa;
    defparam add_17802_6.INJECT1_0 = "NO";
    defparam add_17802_6.INJECT1_1 = "NO";
    CCU2D add_17802_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24462), 
          .COUT(n24463));
    defparam add_17802_4.INIT0 = 16'h5555;
    defparam add_17802_4.INIT1 = 16'h5aaa;
    defparam add_17802_4.INJECT1_0 = "NO";
    defparam add_17802_4.INJECT1_1 = "NO";
    CCU2D add_17802_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24462));
    defparam add_17802_2.INIT0 = 16'h1000;
    defparam add_17802_2.INIT1 = 16'h5555;
    defparam add_17802_2.INJECT1_0 = "NO";
    defparam add_17802_2.INJECT1_1 = "NO";
    FD1S3IX count_2379__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i1.GSR = "ENABLED";
    FD1S3IX count_2379__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i2.GSR = "ENABLED";
    FD1S3IX count_2379__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i3.GSR = "ENABLED";
    FD1S3IX count_2379__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i4.GSR = "ENABLED";
    FD1S3IX count_2379__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i5.GSR = "ENABLED";
    FD1S3IX count_2379__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i6.GSR = "ENABLED";
    FD1S3IX count_2379__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i7.GSR = "ENABLED";
    FD1S3IX count_2379__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i8.GSR = "ENABLED";
    FD1S3IX count_2379__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i9.GSR = "ENABLED";
    FD1S3IX count_2379__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i10.GSR = "ENABLED";
    FD1S3IX count_2379__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i11.GSR = "ENABLED";
    FD1S3IX count_2379__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i12.GSR = "ENABLED";
    FD1S3IX count_2379__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i13.GSR = "ENABLED";
    FD1S3IX count_2379__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i14.GSR = "ENABLED";
    FD1S3IX count_2379__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i15.GSR = "ENABLED";
    FD1S3IX count_2379__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i16.GSR = "ENABLED";
    FD1S3IX count_2379__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i17.GSR = "ENABLED";
    FD1S3IX count_2379__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i18.GSR = "ENABLED";
    FD1S3IX count_2379__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i19.GSR = "ENABLED";
    FD1S3IX count_2379__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i20.GSR = "ENABLED";
    FD1S3IX count_2379__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i21.GSR = "ENABLED";
    FD1S3IX count_2379__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i22.GSR = "ENABLED";
    FD1S3IX count_2379__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i23.GSR = "ENABLED";
    FD1S3IX count_2379__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i24.GSR = "ENABLED";
    FD1S3IX count_2379__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i25.GSR = "ENABLED";
    FD1S3IX count_2379__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i26.GSR = "ENABLED";
    FD1S3IX count_2379__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i27.GSR = "ENABLED";
    FD1S3IX count_2379__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i28.GSR = "ENABLED";
    FD1S3IX count_2379__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i29.GSR = "ENABLED";
    FD1S3IX count_2379__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i30.GSR = "ENABLED";
    FD1S3IX count_2379__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n14872), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2379__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000) 
//

module \ClockDividerP(factor=12000)  (GND_net, debug_c_c, n2736, select_clk, 
            n16717, n7591, n28406, \state[0] , n28477, n28404, n26896) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n2736;
    output select_clk;
    input n16717;
    output n7591;
    output n28406;
    input \state[0] ;
    input n28477;
    output n28404;
    output n26896;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24376;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n24375, n24374, n24373, n24372, n24371, n24370, n24369, 
        n24368, n24367, n24366, n24365, n24364, n24363, n24362, 
        n24361, n24461, n24460, n24459, n24458, n24457, n24456, 
        n24455, n24454, n24453, n24452, n24992, n15, n20, n16, 
        n24451, n27, n40, n36, n28, n18, n38, n32, n24450, 
        n24449, n34, n24;
    
    CCU2D count_2378_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24376), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_33.INIT1 = 16'h0000;
    defparam count_2378_add_4_33.INJECT1_0 = "NO";
    defparam count_2378_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24375), .COUT(n24376), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_31.INJECT1_0 = "NO";
    defparam count_2378_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24374), .COUT(n24375), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_29.INJECT1_0 = "NO";
    defparam count_2378_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24373), .COUT(n24374), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_27.INJECT1_0 = "NO";
    defparam count_2378_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24372), .COUT(n24373), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_25.INJECT1_0 = "NO";
    defparam count_2378_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24371), .COUT(n24372), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_23.INJECT1_0 = "NO";
    defparam count_2378_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24370), .COUT(n24371), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_21.INJECT1_0 = "NO";
    defparam count_2378_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24369), .COUT(n24370), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_19.INJECT1_0 = "NO";
    defparam count_2378_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24368), .COUT(n24369), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_17.INJECT1_0 = "NO";
    defparam count_2378_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24367), .COUT(n24368), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_15.INJECT1_0 = "NO";
    defparam count_2378_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24366), .COUT(n24367), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_13.INJECT1_0 = "NO";
    defparam count_2378_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24365), .COUT(n24366), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_11.INJECT1_0 = "NO";
    defparam count_2378_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24364), .COUT(n24365), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_9.INJECT1_0 = "NO";
    defparam count_2378_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24363), .COUT(n24364), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_7.INJECT1_0 = "NO";
    defparam count_2378_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24362), .COUT(n24363), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_5.INJECT1_0 = "NO";
    defparam count_2378_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24361), .COUT(n24362), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2378_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2378_add_4_3.INJECT1_0 = "NO";
    defparam count_2378_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2378_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24361), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378_add_4_1.INIT0 = 16'hF000;
    defparam count_2378_add_4_1.INIT1 = 16'h0555;
    defparam count_2378_add_4_1.INJECT1_0 = "NO";
    defparam count_2378_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2378__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2736), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i0.GSR = "ENABLED";
    FD1S3AX clk_o_14 (.D(n16717), .CK(debug_c_c), .Q(select_clk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=25, LSE_RCOL=48, LSE_LLINE=21, LSE_RLINE=23 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_285 (.A(n7591), .B(select_clk), .Z(n28406)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam i1_2_lut_rep_285.init = 16'h2222;
    FD1S3IX count_2378__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2736), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i1.GSR = "ENABLED";
    CCU2D add_17803_28 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24461), 
          .S1(n7591));
    defparam add_17803_28.INIT0 = 16'h5555;
    defparam add_17803_28.INIT1 = 16'h0000;
    defparam add_17803_28.INJECT1_0 = "NO";
    defparam add_17803_28.INJECT1_1 = "NO";
    CCU2D add_17803_26 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24460), .COUT(n24461));
    defparam add_17803_26.INIT0 = 16'h5555;
    defparam add_17803_26.INIT1 = 16'h5555;
    defparam add_17803_26.INJECT1_0 = "NO";
    defparam add_17803_26.INJECT1_1 = "NO";
    CCU2D add_17803_24 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24459), .COUT(n24460));
    defparam add_17803_24.INIT0 = 16'h5555;
    defparam add_17803_24.INIT1 = 16'h5555;
    defparam add_17803_24.INJECT1_0 = "NO";
    defparam add_17803_24.INJECT1_1 = "NO";
    CCU2D add_17803_22 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24458), .COUT(n24459));
    defparam add_17803_22.INIT0 = 16'h5555;
    defparam add_17803_22.INIT1 = 16'h5555;
    defparam add_17803_22.INJECT1_0 = "NO";
    defparam add_17803_22.INJECT1_1 = "NO";
    CCU2D add_17803_20 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24457), .COUT(n24458));
    defparam add_17803_20.INIT0 = 16'h5555;
    defparam add_17803_20.INIT1 = 16'h5555;
    defparam add_17803_20.INJECT1_0 = "NO";
    defparam add_17803_20.INJECT1_1 = "NO";
    CCU2D add_17803_18 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24456), .COUT(n24457));
    defparam add_17803_18.INIT0 = 16'h5555;
    defparam add_17803_18.INIT1 = 16'h5555;
    defparam add_17803_18.INJECT1_0 = "NO";
    defparam add_17803_18.INJECT1_1 = "NO";
    CCU2D add_17803_16 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24455), .COUT(n24456));
    defparam add_17803_16.INIT0 = 16'h5555;
    defparam add_17803_16.INIT1 = 16'h5555;
    defparam add_17803_16.INJECT1_0 = "NO";
    defparam add_17803_16.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_283_4_lut (.A(n7591), .B(select_clk), .C(\state[0] ), 
         .D(n28477), .Z(n28404)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam i1_3_lut_rep_283_4_lut.init = 16'h0002;
    FD1S3IX count_2378__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2736), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i2.GSR = "ENABLED";
    FD1S3IX count_2378__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2736), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i3.GSR = "ENABLED";
    FD1S3IX count_2378__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2736), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i4.GSR = "ENABLED";
    FD1S3IX count_2378__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2736), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i5.GSR = "ENABLED";
    FD1S3IX count_2378__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2736), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i6.GSR = "ENABLED";
    FD1S3IX count_2378__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2736), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i7.GSR = "ENABLED";
    FD1S3IX count_2378__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2736), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i8.GSR = "ENABLED";
    FD1S3IX count_2378__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2736), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i9.GSR = "ENABLED";
    FD1S3IX count_2378__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i10.GSR = "ENABLED";
    FD1S3IX count_2378__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i11.GSR = "ENABLED";
    FD1S3IX count_2378__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i12.GSR = "ENABLED";
    FD1S3IX count_2378__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i13.GSR = "ENABLED";
    FD1S3IX count_2378__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i14.GSR = "ENABLED";
    FD1S3IX count_2378__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i15.GSR = "ENABLED";
    FD1S3IX count_2378__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i16.GSR = "ENABLED";
    FD1S3IX count_2378__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i17.GSR = "ENABLED";
    FD1S3IX count_2378__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i18.GSR = "ENABLED";
    FD1S3IX count_2378__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i19.GSR = "ENABLED";
    FD1S3IX count_2378__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i20.GSR = "ENABLED";
    FD1S3IX count_2378__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i21.GSR = "ENABLED";
    FD1S3IX count_2378__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i22.GSR = "ENABLED";
    FD1S3IX count_2378__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i23.GSR = "ENABLED";
    FD1S3IX count_2378__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i24.GSR = "ENABLED";
    FD1S3IX count_2378__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i25.GSR = "ENABLED";
    FD1S3IX count_2378__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i26.GSR = "ENABLED";
    FD1S3IX count_2378__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i27.GSR = "ENABLED";
    FD1S3IX count_2378__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i28.GSR = "ENABLED";
    FD1S3IX count_2378__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i29.GSR = "ENABLED";
    FD1S3IX count_2378__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i30.GSR = "ENABLED";
    FD1S3IX count_2378__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2736), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2378__i31.GSR = "ENABLED";
    CCU2D add_17803_14 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24454), .COUT(n24455));
    defparam add_17803_14.INIT0 = 16'h5555;
    defparam add_17803_14.INIT1 = 16'h5555;
    defparam add_17803_14.INJECT1_0 = "NO";
    defparam add_17803_14.INJECT1_1 = "NO";
    CCU2D add_17803_12 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24453), .COUT(n24454));
    defparam add_17803_12.INIT0 = 16'h5555;
    defparam add_17803_12.INIT1 = 16'h5555;
    defparam add_17803_12.INJECT1_0 = "NO";
    defparam add_17803_12.INJECT1_1 = "NO";
    CCU2D add_17803_10 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24452), .COUT(n24453));
    defparam add_17803_10.INIT0 = 16'h5555;
    defparam add_17803_10.INIT1 = 16'h5555;
    defparam add_17803_10.INJECT1_0 = "NO";
    defparam add_17803_10.INJECT1_1 = "NO";
    LUT4 i20297_4_lut (.A(n24992), .B(n15), .C(n20), .D(n16), .Z(n26896)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i20297_4_lut.init = 16'h4000;
    CCU2D add_17803_8 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24451), .COUT(n24452));
    defparam add_17803_8.INIT0 = 16'h5555;
    defparam add_17803_8.INIT1 = 16'h5aaa;
    defparam add_17803_8.INJECT1_0 = "NO";
    defparam add_17803_8.INJECT1_1 = "NO";
    LUT4 i20_4_lut (.A(n27), .B(n40), .C(n36), .D(n28), .Z(n24992)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[11]), .B(count[10]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(count[9]), .B(n18), .C(count[6]), .D(count[7]), 
         .Z(n20)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(count[1]), .B(count[4]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i6_2_lut (.A(count[28]), .B(count[12]), .Z(n27)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[5]), .B(n38), .C(n32), .D(count[20]), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(count[8]), .B(count[25]), .C(count[15]), .D(count[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[17]), .B(count[24]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i7_4_lut (.A(count[13]), .B(count[2]), .C(count[3]), .D(count[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    CCU2D add_17803_6 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24450), .COUT(n24451));
    defparam add_17803_6.INIT0 = 16'h5aaa;
    defparam add_17803_6.INIT1 = 16'h5aaa;
    defparam add_17803_6.INJECT1_0 = "NO";
    defparam add_17803_6.INJECT1_1 = "NO";
    CCU2D add_17803_4 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24449), 
          .COUT(n24450));
    defparam add_17803_4.INIT0 = 16'h5555;
    defparam add_17803_4.INIT1 = 16'h5aaa;
    defparam add_17803_4.INJECT1_0 = "NO";
    defparam add_17803_4.INJECT1_1 = "NO";
    CCU2D add_17803_2 (.A0(count[5]), .B0(count[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24449));
    defparam add_17803_2.INIT0 = 16'h7000;
    defparam add_17803_2.INIT1 = 16'h5aaa;
    defparam add_17803_2.INJECT1_0 = "NO";
    defparam add_17803_2.INJECT1_1 = "NO";
    LUT4 i17_4_lut (.A(count[29]), .B(n34), .C(n24), .D(count[14]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(count[22]), .B(count[21]), .C(count[31]), .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(count[16]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[19]), .B(count[18]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (register_addr, n11, n12585, n26425, 
            n19316, rw, n28415, debug_c_c, n30473, n28485, databus_out, 
            \select[7] , debug_c_2, \select[2] , n28457, \select[1] , 
            n28542, n28438, n26396, n28441, prev_select, n28477, 
            n3539, \sendcount[1] , n30468, databus, \read_value[5] , 
            n4, \read_value[7] , n4_adj_147, \read_value[0] , n4_adj_148, 
            \read_value[3] , n4_adj_149, \read_value[2] , n4_adj_150, 
            \read_value[4] , n4_adj_151, n8, \read_size[0] , \read_value[6] , 
            n4_adj_152, n52, \read_value[13] , n2, \read_value[10] , 
            n2_adj_153, \read_value[26] , n2_adj_154, \read_value[31] , 
            n2_adj_155, \read_value[29] , n2_adj_156, \read_value[9] , 
            n2_adj_157, \read_value[11] , n2_adj_158, \read_value[30] , 
            n2_adj_159, \read_value[28] , n2_adj_160, \read_value[27] , 
            n2_adj_161, \read_value[25] , n2_adj_162, \read_value[24] , 
            n2_adj_163, \read_value[23] , n2_adj_164, \read_value[22] , 
            n2_adj_165, \read_value[21] , n2_adj_166, \read_value[20] , 
            n2_adj_167, \read_value[19] , n2_adj_168, \read_value[18] , 
            n2_adj_169, \read_value[17] , n2_adj_170, \read_value[16] , 
            n2_adj_171, \read_value[15] , n2_adj_172, \read_value[14] , 
            n2_adj_173, \read_value[12] , n2_adj_174, n11943, n28563, 
            \read_value[8] , n2_adj_175, n28442, n9, n10, debug_c_7, 
            \reg_size[2] , n28576, n28431, prev_select_adj_176, n28414, 
            n28482, n151, n12649, n28430, n3356, prev_select_adj_177, 
            n30467, \read_value[23]_adj_178 , n1, \read_value[22]_adj_179 , 
            n1_adj_180, n26540, n8273, n3452, debug_c_3, \register[2][14] , 
            n26079, \register[2][12] , n26098, \register[2][10] , n26081, 
            \register[2][7] , n26090, \register[2][11] , n26083, n28448, 
            n28452, \control_reg[7] , n7685, \control_reg[7]_adj_181 , 
            n7694, \register[2][6] , n26088, \register[2][5] , n26096, 
            \register[2][9] , n26077, \register[2][8] , n26076, \register[2][13] , 
            n26085, \register[2][4] , n26100, n28440, n14798, n26514, 
            \register[2][15] , n26087, \control_reg[7]_adj_182 , n7703, 
            n28451, \register[2][16] , n26084, \register[2][17] , n26094, 
            \register[2][18] , n26095, \steps_reg[5] , n14, \register[2][19] , 
            n26093, \register[2][20] , n26091, \register[2][21] , n26092, 
            \read_value[21]_adj_183 , n1_adj_184, n28480, \register[2][22] , 
            n26080, \register[2][23] , n26086, n28458, \register[2][24] , 
            n26078, \register[2][25] , n26082, \register[2][26] , n26089, 
            \register[2][27] , n26102, \register[2][28] , n26097, \register[2][29] , 
            n26099, \register[2][30] , n26103, n3626, n26489, n28476, 
            n28487, n26437, n26439, n233, \register[2][31] , n26101, 
            prev_select_adj_185, n8472, \steps_reg[6] , n13, \steps_reg[3] , 
            n12, \read_value[20]_adj_186 , n1_adj_187, debug_c_4, \read_value[19]_adj_188 , 
            n1_adj_189, \read_value[18]_adj_190 , n1_adj_191, \read_value[17]_adj_192 , 
            n1_adj_193, n12981, \read_value[16]_adj_194 , n1_adj_195, 
            n15, n8336, n4_adj_196, n12580, n62, n15_adj_197, n27504, 
            n27505, n27502, n27503, n28425, n28439, n176, \read_value[15]_adj_198 , 
            n1_adj_199, debug_c_5, \read_value[14]_adj_200 , n1_adj_201, 
            \read_value[12]_adj_202 , n1_adj_203, \read_value[8]_adj_204 , 
            n1_adj_205, n12647, \read_value[10]_adj_206 , n1_adj_207, 
            \read_value[30]_adj_208 , n1_adj_209, n12599, \read_value[9]_adj_210 , 
            n1_adj_211, \read_value[11]_adj_212 , n1_adj_213, \read_value[13]_adj_214 , 
            n1_adj_215, n28445, \read_value[27]_adj_216 , n1_adj_217, 
            \read_value[28]_adj_218 , n1_adj_219, \read_value[31]_adj_220 , 
            n1_adj_221, \read_value[29]_adj_222 , n1_adj_223, \read_value[1] , 
            n1_adj_224, \read_value[26]_adj_225 , n1_adj_226, n12995, 
            \read_value[25]_adj_227 , n1_adj_228, \read_value[24]_adj_229 , 
            n1_adj_230, \steps_reg[7] , n12_adj_231, \reset_count[7] , 
            \reset_count[6] , \reset_count[5] , n24551, n9969, GND_net, 
            n9970_c) /* synthesis syn_module_defined=1 */ ;
    output [7:0]register_addr;
    input n11;
    input n12585;
    output n26425;
    output n19316;
    output rw;
    output n28415;
    input debug_c_c;
    input n30473;
    input n28485;
    output [31:0]databus_out;
    output \select[7] ;
    output debug_c_2;
    output \select[2] ;
    input n28457;
    output \select[1] ;
    output n28542;
    output n28438;
    output n26396;
    output n28441;
    input prev_select;
    input n28477;
    output n3539;
    output \sendcount[1] ;
    output n30468;
    input [31:0]databus;
    input \read_value[5] ;
    output n4;
    input \read_value[7] ;
    output n4_adj_147;
    input \read_value[0] ;
    output n4_adj_148;
    input \read_value[3] ;
    output n4_adj_149;
    input \read_value[2] ;
    output n4_adj_150;
    input \read_value[4] ;
    output n4_adj_151;
    input n8;
    input \read_size[0] ;
    input \read_value[6] ;
    output n4_adj_152;
    output n52;
    input \read_value[13] ;
    output n2;
    input \read_value[10] ;
    output n2_adj_153;
    input \read_value[26] ;
    output n2_adj_154;
    input \read_value[31] ;
    output n2_adj_155;
    input \read_value[29] ;
    output n2_adj_156;
    input \read_value[9] ;
    output n2_adj_157;
    input \read_value[11] ;
    output n2_adj_158;
    input \read_value[30] ;
    output n2_adj_159;
    input \read_value[28] ;
    output n2_adj_160;
    input \read_value[27] ;
    output n2_adj_161;
    input \read_value[25] ;
    output n2_adj_162;
    input \read_value[24] ;
    output n2_adj_163;
    input \read_value[23] ;
    output n2_adj_164;
    input \read_value[22] ;
    output n2_adj_165;
    input \read_value[21] ;
    output n2_adj_166;
    input \read_value[20] ;
    output n2_adj_167;
    input \read_value[19] ;
    output n2_adj_168;
    input \read_value[18] ;
    output n2_adj_169;
    input \read_value[17] ;
    output n2_adj_170;
    input \read_value[16] ;
    output n2_adj_171;
    input \read_value[15] ;
    output n2_adj_172;
    input \read_value[14] ;
    output n2_adj_173;
    input \read_value[12] ;
    output n2_adj_174;
    input n11943;
    output n28563;
    input \read_value[8] ;
    output n2_adj_175;
    output n28442;
    input n9;
    input n10;
    output debug_c_7;
    input \reg_size[2] ;
    input n28576;
    output n28431;
    input prev_select_adj_176;
    output n28414;
    output n28482;
    output n151;
    output n12649;
    input n28430;
    output n3356;
    input prev_select_adj_177;
    input n30467;
    input \read_value[23]_adj_178 ;
    output n1;
    input \read_value[22]_adj_179 ;
    output n1_adj_180;
    output n26540;
    output n8273;
    output n3452;
    output debug_c_3;
    input \register[2][14] ;
    output n26079;
    input \register[2][12] ;
    output n26098;
    input \register[2][10] ;
    output n26081;
    input \register[2][7] ;
    output n26090;
    input \register[2][11] ;
    output n26083;
    output n28448;
    output n28452;
    input \control_reg[7] ;
    output n7685;
    input \control_reg[7]_adj_181 ;
    output n7694;
    input \register[2][6] ;
    output n26088;
    input \register[2][5] ;
    output n26096;
    input \register[2][9] ;
    output n26077;
    input \register[2][8] ;
    output n26076;
    input \register[2][13] ;
    output n26085;
    input \register[2][4] ;
    output n26100;
    output n28440;
    output n14798;
    output n26514;
    input \register[2][15] ;
    output n26087;
    input \control_reg[7]_adj_182 ;
    output n7703;
    output n28451;
    input \register[2][16] ;
    output n26084;
    input \register[2][17] ;
    output n26094;
    input \register[2][18] ;
    output n26095;
    input \steps_reg[5] ;
    output n14;
    input \register[2][19] ;
    output n26093;
    input \register[2][20] ;
    output n26091;
    input \register[2][21] ;
    output n26092;
    input \read_value[21]_adj_183 ;
    output n1_adj_184;
    output n28480;
    input \register[2][22] ;
    output n26080;
    input \register[2][23] ;
    output n26086;
    output n28458;
    input \register[2][24] ;
    output n26078;
    input \register[2][25] ;
    output n26082;
    input \register[2][26] ;
    output n26089;
    input \register[2][27] ;
    output n26102;
    input \register[2][28] ;
    output n26097;
    input \register[2][29] ;
    output n26099;
    input \register[2][30] ;
    output n26103;
    output n3626;
    output n26489;
    output n28476;
    output n28487;
    output n26437;
    output n26439;
    output n233;
    input \register[2][31] ;
    output n26101;
    input prev_select_adj_185;
    output n8472;
    input \steps_reg[6] ;
    output n13;
    input \steps_reg[3] ;
    output n12;
    input \read_value[20]_adj_186 ;
    output n1_adj_187;
    output debug_c_4;
    input \read_value[19]_adj_188 ;
    output n1_adj_189;
    input \read_value[18]_adj_190 ;
    output n1_adj_191;
    input \read_value[17]_adj_192 ;
    output n1_adj_193;
    output n12981;
    input \read_value[16]_adj_194 ;
    output n1_adj_195;
    output n15;
    output n8336;
    output n4_adj_196;
    output n12580;
    output n62;
    output n15_adj_197;
    input n27504;
    output n27505;
    input n27502;
    output n27503;
    output n28425;
    output n28439;
    output n176;
    input \read_value[15]_adj_198 ;
    output n1_adj_199;
    output debug_c_5;
    input \read_value[14]_adj_200 ;
    output n1_adj_201;
    input \read_value[12]_adj_202 ;
    output n1_adj_203;
    input \read_value[8]_adj_204 ;
    output n1_adj_205;
    output n12647;
    input \read_value[10]_adj_206 ;
    output n1_adj_207;
    input \read_value[30]_adj_208 ;
    output n1_adj_209;
    output n12599;
    input \read_value[9]_adj_210 ;
    output n1_adj_211;
    input \read_value[11]_adj_212 ;
    output n1_adj_213;
    input \read_value[13]_adj_214 ;
    output n1_adj_215;
    output n28445;
    input \read_value[27]_adj_216 ;
    output n1_adj_217;
    input \read_value[28]_adj_218 ;
    output n1_adj_219;
    input \read_value[31]_adj_220 ;
    output n1_adj_221;
    input \read_value[29]_adj_222 ;
    output n1_adj_223;
    input \read_value[1] ;
    output n1_adj_224;
    input \read_value[26]_adj_225 ;
    output n1_adj_226;
    output n12995;
    input \read_value[25]_adj_227 ;
    output n1_adj_228;
    input \read_value[24]_adj_229 ;
    output n1_adj_230;
    input \steps_reg[7] ;
    output n12_adj_231;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n24551;
    output n9969;
    input GND_net;
    input n9970_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire n30467 /* synthesis nomerge= */ ;
    
    wire n28459, n2537;
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    wire [31:0]n1278;
    wire [7:0]n2020;
    
    wire n10_c, n26788, n30;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n4_c;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n13149, n25671;
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n26570, n26569, n28455;
    wire [4:0]n18;
    wire [3:0]n8521;
    
    wire n2592;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n28534, n26631, n2594;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n28449, n14664, n12642, n27982;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n28535, n5020, n14803, n28536, n9_c;
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n4_adj_300, n12544, n6, n28486, n26360, n14666;
    wire [127:0]select;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    
    wire n14670, n4_adj_301, n8_c, n14662, n14678;
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]n5011;
    
    wire n28594, n30464, n14676;
    wire [7:0]register_addr_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire n4_adj_302, n28547, n28466, n26399, n28475;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n12174, n14807, n28500, n28428, n27815, n28468;
    wire [4:0]n19;
    
    wire n28517, n28578, n28474, n28548, n28587, n28497, n5, n24767, 
        n26454, n26389, n24764, n28586, n28593, n28592, n24770, 
        n24760, n24771, n24761, n8417, n24756, n24776, n24775, 
        n24762, n24777, n24782, n24753, n24763, n24781, n24797, 
        n24757, n24796, n24800, n24802, n24653, n24798, n24654, 
        n24783, n24656, n24658, n24780, n24660, n24661, n24659, 
        n24662, n28596, n24808, n25655, n25679, n28595, n25677, 
        n25657, n28599, n25741, n25729, n25743, n25693, n25695, 
        n25651, n25727, n28598, n25659, n25681, n25675, n25673, 
        n14669, n14661, n5_adj_305, n28602, n14665, n28601, escape, 
        n9903, n14677, n28605, n28604, n28608, n28607, n29188, 
        n29190, n28611, n28610, n28614, n28613, n11_adj_306, n14_c, 
        n5_adj_307, n26387, n28514, n5_adj_309, n26386, n28583, 
        n4_adj_311, n5_adj_313, n26385, n27976, n11_adj_318, n5_adj_320, 
        n26384, n28584, n5_adj_321, n26383, n28510, n5_adj_322, 
        n26382, n5_adj_323, n26381, n7, n26724, n28579, n5_adj_324, 
        n26380, n1679, n28519, n5_adj_327, n26379, n5_adj_342, n26372, 
        n5_adj_346, n26378, n5_adj_349, n26377, n5_adj_350, n26376, 
        n1_c, n6_adj_352, n9_adj_353, n5_adj_354, n26375, n26578, 
        n28564, n27600, n27601, n26403, n28565, n28481, n28496, 
        n12374, n1383, n5_adj_359, n26371, n5_adj_360, n26373, n28567, 
        n5_adj_361, n26374, n5_adj_362, n26370, n28566, n5_adj_363, 
        n26369, n28511, n5_adj_364, n26368, n28447, n28509;
    wire [3:0]n1674;
    
    wire n28574, n4_adj_365, n28609;
    wire [7:0]n9241;
    
    wire n5_adj_366, n26359, n4_adj_367, n28606, n4_adj_368, n28600, 
        n28577, n26464, n14675, n5_adj_369, n26358, n26579, n26363, 
        n183, n26183, n26298, n14663, n24846, send, n2029, n24779, 
        n5_adj_371, n26367, n5_adj_372, n26366, n27980, n12_c, n26552, 
        n26553, n28518, n27797, n1731, n24909, n24969, n11426, 
        n5_adj_377, n26365, n5_adj_378, n26364, n28580, n8_adj_379, 
        n28585, n5_adj_380, n26362, n5_adj_381, n26361, n28588, 
        n28597, n28603, n5_adj_383, n26388, n28615, n27981, n11_adj_384, 
        n11_adj_385, n11_adj_386, n11_adj_387, n11_adj_388, n11_adj_389, 
        n26299, n25771, n11_adj_390, n11_adj_391, n11_adj_393, n11252, 
        n15_c, n26738, n11_adj_395, n10029, n25785, n11254, n10023, 
        n1390, n1389, n11_adj_398, n25885, n12121, n11_adj_399, 
        n11_adj_400, n11_adj_401, n11_adj_402, n6_adj_403, n28419, 
        n8_adj_404, n8_adj_423, n27814, n5_adj_434, busy, n38, n8_adj_452, 
        n35, n55, n26319, n6_adj_458, n28581;
    
    LUT4 i1_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(n28459), .C(n11), 
         .D(n12585), .Z(n26425)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 mux_500_i1_3_lut (.A(n2537), .B(esc_data[0]), .C(n1278[18]), 
         .Z(n2020[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_500_i1_3_lut.init = 16'hcaca;
    LUT4 i20358_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(n28459), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n19316)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i20358_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i19988_2_lut_rep_294_3_lut_4_lut (.A(register_addr[2]), .B(n28459), 
         .C(rw), .D(register_addr[1]), .Z(n28415)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19988_2_lut_rep_294_3_lut_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut (.A(esc_data[0]), .B(n10_c), .C(n26788), .D(n30), 
         .Z(n2537)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_4_lut.init = 16'h8808;
    LUT4 i4_4_lut (.A(n1278[15]), .B(esc_data[6]), .C(esc_data[5]), .D(esc_data[7]), 
         .Z(n10_c)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut.init = 16'h0002;
    LUT4 i20094_4_lut (.A(esc_data[2]), .B(esc_data[1]), .C(esc_data[4]), 
         .D(esc_data[3]), .Z(n26788)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20094_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(esc_data[4]), .B(esc_data[2]), .C(esc_data[1]), 
         .D(esc_data[3]), .Z(n30)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'h2080;
    LUT4 i1_2_lut (.A(sendcount[0]), .B(sendcount[3]), .Z(n4_c)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut.init = 16'h4444;
    FD1P3IX buffer_0___i1 (.D(n25671), .SP(n13149), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n26570)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_199 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n26569)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_199.init = 16'hfbfb;
    FD1P3AX sendcount__i0 (.D(n18[0]), .SP(n28455), .CK(debug_c_c), .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    LUT4 i13031_2_lut (.A(sendcount[3]), .B(sendcount[0]), .Z(n8521[0])) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i13031_2_lut.init = 16'hdddd;
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    LUT4 i4_2_lut_rep_413 (.A(n1278[14]), .B(n1278[15]), .Z(n28534)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_413.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_200 (.A(n1278[14]), .B(n1278[15]), .C(n1278[12]), 
         .Z(n26631)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_200.init = 16'hfefe;
    LUT4 i918_2_lut (.A(n1278[5]), .B(n28485), .Z(n2594)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i918_2_lut.init = 16'h8888;
    FD1P3AX tx_data_i0_i0 (.D(n2020[0]), .SP(n28449), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n14664), .CK(debug_c_c), .CD(n30473), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n27982), .SP(n12642), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_414 (.A(n1278[19]), .B(n1278[3]), .C(n1278[11]), 
         .Z(n28535)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_rep_414.init = 16'hfefe;
    LUT4 i1_4_lut_adj_201 (.A(n5020), .B(n8521[0]), .C(n28485), .D(n1278[14]), 
         .Z(n14803)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_201.init = 16'h8000;
    LUT4 i3_2_lut_4_lut (.A(n1278[19]), .B(n1278[3]), .C(n1278[11]), .D(n28536), 
         .Z(n9_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_415 (.A(n1278[7]), .B(n1278[13]), .C(n1278[5]), 
         .Z(n28536)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_rep_415.init = 16'hfefe;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_300)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    FD1S3JX state_FSM_i1 (.D(n12544), .CK(debug_c_c), .PD(n30473), .Q(n1278[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n1278[7]), .B(n1278[13]), .C(n1278[5]), .D(n1278[6]), 
         .Z(n6)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_202 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [6]), 
         .Z(n26360)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_202.init = 16'h2020;
    FD1S3IX select__i7 (.D(n14666), .CK(debug_c_c), .CD(n30473), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    FD1S3IX select__i4 (.D(n14670), .CK(debug_c_c), .CD(n30473), .Q(select[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_301)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 i5_4_lut_adj_203 (.A(n9_c), .B(n1278[15]), .C(n8_c), .D(n1278[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_4_lut_adj_203.init = 16'hfffe;
    FD1S3IX select__i2 (.D(n14662), .CK(debug_c_c), .CD(n28457), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1S3IX select__i1 (.D(n14678), .CK(debug_c_c), .CD(n28457), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2594), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i4 (.D(n5011[4]), .SP(n12642), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n5011[2]), .SP(n12642), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n5011[1]), .SP(n12642), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    FD1S3IX bufcount__i3 (.D(n28594), .CK(debug_c_c), .CD(n28457), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n30464), .CK(debug_c_c), .CD(n28457), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n14676), .CK(debug_c_c), .CD(n28457), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2020[4]), .SP(n28449), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2020[3]), .SP(n28449), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2020[1]), .SP(n28449), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr_c[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr_c[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr_c[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2592), .CK(debug_c_c), 
            .Q(register_addr[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_302)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_rep_421 (.A(register_addr[0]), .B(register_addr[1]), .Z(n28542)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_421.init = 16'h4444;
    LUT4 i2_3_lut_rep_317_4_lut (.A(register_addr[0]), .B(register_addr[1]), 
         .C(n28547), .D(n28466), .Z(n28438)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_317_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_320_3_lut (.A(register_addr[0]), .B(register_addr[1]), 
         .C(n26396), .Z(n28441)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_320_3_lut.init = 16'h4040;
    LUT4 i3_4_lut (.A(prev_select), .B(n26399), .C(n28477), .D(n28475), 
         .Z(n3539)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i13932_3_lut_rep_328 (.A(n2537), .B(n28485), .C(n1278[18]), .Z(n28449)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i13932_3_lut_rep_328.init = 16'hc8c8;
    LUT4 i1_2_lut_3_lut_adj_204 (.A(rx_data[1]), .B(rx_data[4]), .C(rx_data[3]), 
         .Z(n12174)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_3_lut_adj_204.init = 16'h0808;
    LUT4 i20314_2_lut_3_lut (.A(n2537), .B(n28485), .C(n1278[18]), .Z(n14807)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i20314_2_lut_3_lut.init = 16'h0808;
    LUT4 i263_2_lut_rep_426 (.A(register_addr[2]), .B(register_addr_c[4]), 
         .Z(n28547)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i263_2_lut_rep_426.init = 16'heeee;
    LUT4 i265_2_lut_rep_379_3_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(register_addr[1]), .Z(n28500)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i265_2_lut_rep_379_3_lut.init = 16'hfefe;
    FD1P3IX sendcount__i4 (.D(n27815), .SP(n28455), .CD(n28428), .CK(debug_c_c), 
            .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 i267_2_lut_rep_347_3_lut_4_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n28468)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i267_2_lut_rep_347_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX sendcount__i3 (.D(n19[3]), .SP(n28455), .CD(n28428), .CK(debug_c_c), 
            .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3IX sendcount__i2 (.D(n19[2]), .SP(n28455), .CD(n28428), .CK(debug_c_c), 
            .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n19[1]), .SP(n28455), .CD(n28428), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_396_3_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(select[4]), .Z(n28517)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_396_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_353_3_lut_4_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(n28578), .D(register_addr_c[5]), .Z(n28474)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_353_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_427 (.A(select[4]), .B(n30468), .Z(n28548)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_427.init = 16'h2222;
    LUT4 i20144_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n28587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20144_then_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_376_3_lut (.A(select[4]), .B(n30468), .C(register_addr_c[5]), 
         .Z(n28497)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_376_3_lut.init = 16'h2020;
    LUT4 i2_4_lut (.A(databus[30]), .B(n5), .C(n1278[13]), .D(n26360), 
         .Z(n24767)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 i2_3_lut_4_lut (.A(select[4]), .B(rw), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n26399)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_205 (.A(select[4]), .B(rw), .C(register_addr_c[5]), 
         .Z(n26454)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_205.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_adj_206 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [5]), 
         .Z(n26389)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_206.init = 16'h2020;
    FD1P3IX buffer_0___i48 (.D(n24764), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 i20144_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n28586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20144_else_3_lut.init = 16'hcaca;
    LUT4 select_1894_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1278[4]), 
         .C(rx_data[6]), .D(n26570), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i8667_then_4_lut (.A(bufcount[3]), .B(n1278[0]), .C(n1278[3]), 
         .D(n1278[4]), .Z(n28593)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8667_then_4_lut.init = 16'haaa2;
    FD1P3IX buffer_0___i47 (.D(n24767), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    LUT4 i8667_else_4_lut (.A(bufcount[3]), .B(n1278[0]), .C(n1278[3]), 
         .D(n1278[4]), .Z(n28592)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8667_else_4_lut.init = 16'h0002;
    FD1P3IX buffer_0___i46 (.D(n24770), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n24760), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n24771), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n24761), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n24756), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n24776), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n24775), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n24762), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n24777), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n24782), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n24753), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n24763), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n24781), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n24797), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n24757), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n24796), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n24800), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n24802), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n24653), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n24798), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n24654), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n24783), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n24656), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i23 (.D(n24658), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i22 (.D(n24780), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n24660), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n24661), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n24659), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n24662), .SP(n13149), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    LUT4 i20147_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n28596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20147_then_3_lut.init = 16'hcaca;
    FD1P3IX buffer_0___i17 (.D(n24808), .SP(n13149), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n25655), .SP(n13149), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n25679), .SP(n13149), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    LUT4 i20147_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n28595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20147_else_3_lut.init = 16'hcaca;
    FD1P3IX buffer_0___i14 (.D(n25677), .SP(n13149), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n25657), .SP(n13149), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    LUT4 i20150_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n28599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20150_then_3_lut.init = 16'hcaca;
    FD1P3IX buffer_0___i12 (.D(n25741), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n25729), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n25743), .SP(n8417), .CD(n28457), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n25693), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n25695), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n25651), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n25727), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    LUT4 i20150_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n28598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20150_else_3_lut.init = 16'hcaca;
    FD1P3IX buffer_0___i5 (.D(n25659), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n25681), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n25675), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i2 (.D(n25673), .SP(n8417), .CD(n30473), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_207 (.A(n1278[0]), .B(n1278[8]), .C(select[4]), 
         .Z(n14669)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_207.init = 16'h1010;
    LUT4 i13108_2_lut_3_lut (.A(n1278[0]), .B(n1278[8]), .C(\select[2] ), 
         .Z(n14661)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i13108_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_4_lut_adj_208 (.A(databus[29]), .B(n5_adj_305), .C(n1278[13]), 
         .D(n26389), .Z(n24770)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_208.init = 16'hffec;
    LUT4 i20153_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n28602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20153_then_3_lut.init = 16'hcaca;
    LUT4 i13158_2_lut_3_lut (.A(n1278[0]), .B(n1278[8]), .C(\select[7] ), 
         .Z(n14665)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i13158_2_lut_3_lut.init = 16'h1010;
    FD1P3AX rw_498 (.D(n1278[10]), .SP(n2592), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i20153_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n28601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20153_else_3_lut.init = 16'hcaca;
    FD1S3AX escape_501 (.D(n9903), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 i13257_2_lut_3_lut (.A(n1278[0]), .B(n1278[8]), .C(\select[1] ), 
         .Z(n14677)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i13257_2_lut_3_lut.init = 16'h1010;
    LUT4 select_1894_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1278[4]), 
         .C(rx_data[5]), .D(n26570), .Z(n5_adj_305)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i20156_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n28605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20156_then_3_lut.init = 16'hcaca;
    LUT4 i20156_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n28604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20156_else_3_lut.init = 16'hcaca;
    LUT4 i20159_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n28608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20159_then_3_lut.init = 16'hcaca;
    LUT4 i20159_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n28607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20159_else_3_lut.init = 16'hcaca;
    LUT4 n29188_bdd_4_lut (.A(n29188), .B(n1278[4]), .C(n29190), .D(bufcount[2]), 
         .Z(n30464)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n29188_bdd_4_lut.init = 16'heef0;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n28611)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n28610)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 i20719_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n28614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20719_then_3_lut.init = 16'hcaca;
    LUT4 i20719_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n28613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20719_else_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_209 (.A(n1278[4]), .B(\buffer[0] [0]), .C(n11_adj_306), 
         .D(n14_c), .Z(n25671)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_209.init = 16'heca0;
    LUT4 i2_4_lut_adj_210 (.A(databus[28]), .B(n5_adj_307), .C(n1278[13]), 
         .D(n26387), .Z(n24760)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_210.init = 16'hffec;
    LUT4 select_1894_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1278[4]), 
         .C(rx_data[4]), .D(n26570), .Z(n5_adj_307)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3956_i4_2_lut_3_lut_4_lut (.A(n28514), .B(n28517), .C(\read_value[5] ), 
         .D(rw), .Z(n4)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3956_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_4_lut_adj_211 (.A(databus[27]), .B(n5_adj_309), .C(n1278[13]), 
         .D(n26386), .Z(n24771)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_211.init = 16'hffec;
    LUT4 Select_3954_i4_2_lut_3_lut_4_lut (.A(n28514), .B(n28517), .C(\read_value[7] ), 
         .D(n30468), .Z(n4_adj_147)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3954_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i20141_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n28583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20141_else_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_311)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 select_1894_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1278[4]), 
         .C(rx_data[3]), .D(n26570), .Z(n5_adj_309)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3961_i4_2_lut_3_lut_4_lut (.A(n28514), .B(n28517), .C(\read_value[0] ), 
         .D(n30468), .Z(n4_adj_148)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3961_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_4_lut_adj_212 (.A(databus[26]), .B(n5_adj_313), .C(n1278[13]), 
         .D(n26385), .Z(n24761)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_212.init = 16'hffec;
    LUT4 select_1894_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1278[4]), 
         .C(rx_data[2]), .D(n26570), .Z(n5_adj_313)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3958_i4_2_lut_3_lut_4_lut (.A(n28514), .B(n28517), .C(\read_value[3] ), 
         .D(rw), .Z(n4_adj_149)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3958_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 n11947_bdd_2_lut_20832 (.A(sendcount[0]), .B(sendcount[3]), .Z(n27976)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n11947_bdd_2_lut_20832.init = 16'hbbbb;
    LUT4 Select_3959_i4_2_lut_3_lut_4_lut (.A(n28514), .B(n28517), .C(\read_value[2] ), 
         .D(n30468), .Z(n4_adj_150)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3959_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3957_i4_2_lut_3_lut_4_lut (.A(n28514), .B(n28517), .C(\read_value[4] ), 
         .D(n30468), .Z(n4_adj_151)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3957_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i4_3_lut_4_lut (.A(n28514), .B(n28517), .C(n8), .D(\read_size[0] ), 
         .Z(n11_adj_318)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4_3_lut_4_lut.init = 16'hf4f0;
    LUT4 Select_3955_i4_2_lut_3_lut_4_lut (.A(n28514), .B(n28517), .C(\read_value[6] ), 
         .D(n30468), .Z(n4_adj_152)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3955_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_4_lut_adj_213 (.A(databus[25]), .B(n5_adj_320), .C(n1278[13]), 
         .D(n26384), .Z(n24756)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_213.init = 16'hffec;
    LUT4 select_1894_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1278[4]), 
         .C(rx_data[1]), .D(n26570), .Z(n5_adj_320)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 i20141_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n28584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20141_then_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_214 (.A(databus[24]), .B(n5_adj_321), .C(n1278[13]), 
         .D(n26383), .Z(n24776)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_214.init = 16'hffec;
    LUT4 select_1894_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1278[4]), 
         .C(rx_data[0]), .D(n26570), .Z(n5_adj_321)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 i20_2_lut_3_lut_4_lut (.A(register_addr_c[5]), .B(n28510), .C(n30468), 
         .D(n28578), .Z(n52)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i20_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i2_4_lut_adj_215 (.A(databus[23]), .B(n5_adj_322), .C(n1278[13]), 
         .D(n26382), .Z(n24775)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_215.init = 16'hffec;
    LUT4 select_1894_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1278[4]), 
         .C(rx_data[7]), .D(n26569), .Z(n5_adj_322)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_216 (.A(databus[22]), .B(n5_adj_323), .C(n1278[13]), 
         .D(n26381), .Z(n24762)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_216.init = 16'hffec;
    LUT4 i20386_4_lut (.A(n7), .B(n26724), .C(n28579), .D(n1278[3]), 
         .Z(n8417)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i20386_4_lut.init = 16'h0544;
    LUT4 select_1894_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1278[4]), 
         .C(rx_data[6]), .D(n26569), .Z(n5_adj_323)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 i20033_3_lut (.A(n1278[13]), .B(n1278[0]), .C(n1278[4]), .Z(n26724)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i20033_3_lut.init = 16'hfefe;
    LUT4 i2_4_lut_adj_217 (.A(databus[21]), .B(n5_adj_324), .C(n1278[13]), 
         .D(n26380), .Z(n24777)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_217.init = 16'hffec;
    LUT4 i486_2_lut (.A(n1278[3]), .B(n1278[4]), .Z(n1679)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i486_2_lut.init = 16'heeee;
    LUT4 select_1894_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1278[4]), 
         .C(rx_data[5]), .D(n26569), .Z(n5_adj_324)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3943_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[13] ), 
         .D(rw), .Z(n2)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3943_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3949_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[10] ), 
         .D(rw), .Z(n2_adj_153)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3949_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3917_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[26] ), 
         .D(rw), .Z(n2_adj_154)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3917_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_218 (.A(databus[20]), .B(n5_adj_327), .C(n1278[13]), 
         .D(n26379), .Z(n24782)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_218.init = 16'hffec;
    LUT4 select_1894_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1278[4]), 
         .C(rx_data[4]), .D(n26569), .Z(n5_adj_327)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3907_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[31] ), 
         .D(rw), .Z(n2_adj_155)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3907_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3911_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[29] ), 
         .D(n30468), .Z(n2_adj_156)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3911_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3951_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[9] ), 
         .D(rw), .Z(n2_adj_157)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3951_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3947_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[11] ), 
         .D(rw), .Z(n2_adj_158)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3947_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3909_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[30] ), 
         .D(rw), .Z(n2_adj_159)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3909_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3913_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[28] ), 
         .D(rw), .Z(n2_adj_160)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3913_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3915_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[27] ), 
         .D(rw), .Z(n2_adj_161)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3915_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3919_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[25] ), 
         .D(rw), .Z(n2_adj_162)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3919_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3921_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[24] ), 
         .D(rw), .Z(n2_adj_163)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3921_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3923_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[23] ), 
         .D(rw), .Z(n2_adj_164)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3923_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3925_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[22] ), 
         .D(rw), .Z(n2_adj_165)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3925_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3927_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[21] ), 
         .D(rw), .Z(n2_adj_166)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3927_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3929_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[20] ), 
         .D(rw), .Z(n2_adj_167)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3929_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3931_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[19] ), 
         .D(rw), .Z(n2_adj_168)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3931_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_219 (.A(databus[19]), .B(n5_adj_342), .C(n1278[13]), 
         .D(n26372), .Z(n24753)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_219.init = 16'hffec;
    LUT4 select_1894_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1278[4]), 
         .C(rx_data[3]), .D(n26569), .Z(n5_adj_342)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3933_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[18] ), 
         .D(rw), .Z(n2_adj_169)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3933_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3935_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[17] ), 
         .D(rw), .Z(n2_adj_170)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3935_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3937_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[16] ), 
         .D(rw), .Z(n2_adj_171)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3937_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_220 (.A(databus[18]), .B(n5_adj_346), .C(n1278[13]), 
         .D(n26378), .Z(n24763)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_220.init = 16'hffec;
    LUT4 select_1894_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1278[4]), 
         .C(rx_data[2]), .D(n26569), .Z(n5_adj_346)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3939_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[15] ), 
         .D(rw), .Z(n2_adj_172)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3939_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3941_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[14] ), 
         .D(rw), .Z(n2_adj_173)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3941_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_221 (.A(databus[17]), .B(n5_adj_349), .C(n1278[13]), 
         .D(n26377), .Z(n24781)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_221.init = 16'hffec;
    LUT4 select_1894_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1278[4]), 
         .C(rx_data[1]), .D(n26569), .Z(n5_adj_349)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_222 (.A(databus[16]), .B(n5_adj_350), .C(n1278[13]), 
         .D(n26376), .Z(n24797)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_222.init = 16'hffec;
    LUT4 Select_3945_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[12] ), 
         .D(rw), .Z(n2_adj_174)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3945_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 select_1894_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1278[4]), 
         .C(rx_data[0]), .D(n26569), .Z(n5_adj_350)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_223 (.A(sendcount[4]), .B(n1_c), .C(n6_adj_352), 
         .D(n11943), .Z(n9_adj_353)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_223.init = 16'hfeff;
    LUT4 i261_2_lut_rep_442 (.A(register_addr[1]), .B(register_addr[0]), 
         .Z(n28563)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i261_2_lut_rep_442.init = 16'heeee;
    LUT4 i2_4_lut_adj_224 (.A(databus[15]), .B(n5_adj_354), .C(n1278[13]), 
         .D(n26375), .Z(n24757)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_224.init = 16'hffec;
    LUT4 Select_3953_i2_2_lut_3_lut_4_lut (.A(n28519), .B(n28517), .C(\read_value[8] ), 
         .D(rw), .Z(n2_adj_175)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3953_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_321_3_lut (.A(register_addr[1]), .B(register_addr[0]), 
         .C(n26396), .Z(n28442)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_321_3_lut.init = 16'h1010;
    LUT4 equal_48_i1_4_lut (.A(sendcount[0]), .B(n11_adj_318), .C(n9), 
         .D(n10), .Z(n1_c)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_48_i1_4_lut.init = 16'h5556;
    LUT4 select_1894_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1278[4]), 
         .C(rx_data[7]), .D(n26578), .Z(n5_adj_354)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_443 (.A(n1278[14]), .B(sendcount[4]), .Z(n28564)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_443.init = 16'h2222;
    LUT4 motor_pwm_r_c_bdd_2_lut_20600_3_lut (.A(n1278[14]), .B(sendcount[4]), 
         .C(n27600), .Z(n27601)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam motor_pwm_r_c_bdd_2_lut_20600_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_adj_225 (.A(n26403), .B(debug_c_7), .C(n1278[0]), .D(n1278[1]), 
         .Z(n12544)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_225.init = 16'hbbba;
    LUT4 i2_4_lut_adj_226 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n28576), .Z(n6_adj_352)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_226.init = 16'he7de;
    LUT4 i1_2_lut_rep_444 (.A(register_addr[2]), .B(register_addr_c[4]), 
         .Z(n28565)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_444.init = 16'h4444;
    LUT4 i1_2_lut_rep_389_3_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(select[4]), .Z(n28510)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_389_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_360_3_lut_4_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(n28578), .D(register_addr_c[5]), .Z(n28481)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_360_3_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_rep_293_4_lut (.A(n28548), .B(n28431), .C(n28542), .D(prev_select_adj_176), 
         .Z(n28414)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_rep_293_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_354_3_lut_4_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(n28578), .D(register_addr_c[5]), .Z(n28475)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_354_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_rep_361_3_lut_4_lut (.A(register_addr[2]), .B(register_addr_c[4]), 
         .C(register_addr_c[5]), .D(select[4]), .Z(n28482)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_361_3_lut_4_lut.init = 16'h0400;
    LUT4 reduce_or_441_i1_3_lut_4_lut (.A(n28496), .B(n12374), .C(\buffer[0] [7]), 
         .D(n1278[9]), .Z(n1383)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_441_i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i2_4_lut_adj_227 (.A(databus[14]), .B(n5_adj_359), .C(n1278[13]), 
         .D(n26371), .Z(n24796)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_227.init = 16'hffec;
    LUT4 select_1894_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1278[4]), 
         .C(rx_data[6]), .D(n26578), .Z(n5_adj_359)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_228 (.A(databus[13]), .B(n5_adj_360), .C(n1278[13]), 
         .D(n26373), .Z(n24800)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_228.init = 16'hffec;
    LUT4 select_1894_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1278[4]), 
         .C(rx_data[5]), .D(n26578), .Z(n5_adj_360)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 i3_4_lut_adj_229 (.A(sendcount[3]), .B(n28567), .C(sendcount[2]), 
         .D(n28564), .Z(n26403)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_229.init = 16'h0200;
    LUT4 i2_4_lut_adj_230 (.A(databus[12]), .B(n5_adj_361), .C(n1278[13]), 
         .D(n26374), .Z(n24802)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_230.init = 16'hffec;
    LUT4 select_1894_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1278[4]), 
         .C(rx_data[4]), .D(n26578), .Z(n5_adj_361)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_231 (.A(databus[11]), .B(n5_adj_362), .C(n1278[13]), 
         .D(n26370), .Z(n24653)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_231.init = 16'hffec;
    LUT4 select_1894_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1278[4]), 
         .C(rx_data[3]), .D(n26578), .Z(n5_adj_362)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i3310_2_lut_rep_445 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n28566)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3310_2_lut_rep_445.init = 16'h8888;
    LUT4 i13930_3_lut_rep_334 (.A(n1278[13]), .B(n28485), .C(n1278[14]), 
         .Z(n28455)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i13930_3_lut_rep_334.init = 16'hc8c8;
    LUT4 i13165_3_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(n9_adj_353), 
         .D(sendcount[2]), .Z(n19[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;
    defparam i13165_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i3313_2_lut_rep_446 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n28567)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3313_2_lut_rep_446.init = 16'heeee;
    LUT4 i20307_2_lut_rep_307_3_lut (.A(n1278[13]), .B(n28485), .C(n1278[14]), 
         .Z(n28428)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i20307_2_lut_rep_307_3_lut.init = 16'h0808;
    LUT4 i2_4_lut_adj_232 (.A(databus[10]), .B(n5_adj_363), .C(n1278[13]), 
         .D(n26369), .Z(n24798)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_232.init = 16'hffec;
    LUT4 select_1894_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1278[4]), 
         .C(rx_data[2]), .D(n26578), .Z(n5_adj_363)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_390_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n28511)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_390_3_lut.init = 16'h1e1e;
    LUT4 i2_4_lut_adj_233 (.A(databus[9]), .B(n5_adj_364), .C(n1278[13]), 
         .D(n26368), .Z(n24654)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_233.init = 16'hffec;
    LUT4 select_1894_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1278[4]), 
         .C(rx_data[1]), .D(n26578), .Z(n5_adj_364)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i3027_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n28447), .C(n28509), 
         .D(bufcount[0]), .Z(n1674[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3027_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n28574), .B(n28511), .C(n4_adj_365), 
         .D(n28609), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i2_4_lut_adj_234 (.A(databus[8]), .B(n5_adj_366), .C(n1278[13]), 
         .D(n26359), .Z(n24783)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_234.init = 16'hffec;
    LUT4 select_1894_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1278[4]), 
         .C(rx_data[0]), .D(n26578), .Z(n5_adj_366)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 i3_4_lut_adj_235 (.A(n151), .B(n28565), .C(n28563), .D(n26454), 
         .Z(n12649)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_4_lut_adj_235.init = 16'h0400;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n28574), .B(n28511), .C(n4_adj_367), 
         .D(n28606), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n28574), .B(n28511), .C(n4_adj_368), 
         .D(n28600), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_adj_236 (.A(n1278[3]), .B(n28486), .C(n1278[13]), 
         .Z(n14_c)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_236.init = 16'hf2f2;
    LUT4 i1_2_lut_3_lut_4_lut_adj_237 (.A(n28577), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n12374), .Z(n26464)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_237.init = 16'h0e00;
    PFUMX i8671 (.BLUT(n14675), .ALUT(n1674[1]), .C0(n1679), .Z(n14676));
    LUT4 i2_4_lut_adj_238 (.A(databus[7]), .B(n5_adj_369), .C(n1278[13]), 
         .D(n26358), .Z(n24656)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_238.init = 16'hffec;
    LUT4 select_1894_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1278[4]), 
         .C(rx_data[7]), .D(n26579), .Z(n5_adj_369)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_239 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [7]), 
         .Z(n26363)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_239.init = 16'h2020;
    LUT4 i13300_2_lut (.A(bufcount[1]), .B(n1278[0]), .Z(n14675)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i13300_2_lut.init = 16'h2222;
    LUT4 i3_4_lut_adj_240 (.A(n183), .B(n28481), .C(n28548), .D(n28430), 
         .Z(n3356)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_4_lut_adj_240.init = 16'h8000;
    LUT4 i20391_3_lut (.A(debug_c_7), .B(n26183), .C(n1278[3]), .Z(n26298)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i20391_3_lut.init = 16'h2020;
    LUT4 i1_3_lut_rep_345_4_lut (.A(n28548), .B(register_addr_c[5]), .C(prev_select_adj_177), 
         .D(n28578), .Z(n28466)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i1_3_lut_rep_345_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_adj_241 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [4]), 
         .Z(n26387)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_241.init = 16'h2020;
    PFUMX i8659 (.BLUT(n14663), .ALUT(n24846), .C0(n1679), .Z(n14664));
    FD1P3IX send_491 (.D(n30467), .SP(n2029), .CD(n24779), .CK(debug_c_c), 
            .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_242 (.A(databus[6]), .B(n5_adj_371), .C(n1278[13]), 
         .D(n26367), .Z(n24658)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_242.init = 16'hffec;
    LUT4 select_1894_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1278[4]), 
         .C(rx_data[6]), .D(n26579), .Z(n5_adj_371)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 i3071_2_lut_rep_453 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n28574)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i3071_2_lut_rep_453.init = 16'h9999;
    LUT4 i2_4_lut_adj_243 (.A(databus[5]), .B(n5_adj_372), .C(n1278[13]), 
         .D(n26366), .Z(n24780)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_243.init = 16'hffec;
    LUT4 n11947_bdd_4_lut_20836_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n27980)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n11947_bdd_4_lut_20836_4_lut.init = 16'h6420;
    LUT4 select_1894_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1278[4]), 
         .C(rx_data[5]), .D(n26579), .Z(n5_adj_372)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_244 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [3]), 
         .Z(n26386)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_244.init = 16'h2020;
    LUT4 i20339_3_lut_4_lut (.A(\buffer[0] [1]), .B(n12_c), .C(\buffer[0] [0]), 
         .D(\buffer[0] [2]), .Z(n26552)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i20339_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_245 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [2]), 
         .Z(n26385)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_245.init = 16'h2020;
    LUT4 i20378_3_lut_4_lut (.A(\buffer[0] [1]), .B(n12_c), .C(\buffer[0] [2]), 
         .D(\buffer[0] [0]), .Z(n26553)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i20378_3_lut_4_lut.init = 16'h0010;
    LUT4 i3_4_lut_adj_246 (.A(rx_data[0]), .B(n28518), .C(n27797), .D(escape), 
         .Z(n26183)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_246.init = 16'h0020;
    LUT4 Select_3923_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[23]_adj_178 ), 
         .D(n30468), .Z(n1)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3923_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3925_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[22]_adj_179 ), 
         .D(n30468), .Z(n1_adj_180)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3925_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i13166_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_adj_353), .Z(n19[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i13166_2_lut_2_lut_3_lut.init = 16'h6f6f;
    PFUMX i8665 (.BLUT(n14669), .ALUT(n26553), .C0(n1731), .Z(n14670));
    PFUMX i8673 (.BLUT(n14677), .ALUT(n26552), .C0(n1731), .Z(n14678));
    PFUMX i8661 (.BLUT(n14665), .ALUT(n24909), .C0(n1731), .Z(n14666));
    PFUMX i8657 (.BLUT(n14661), .ALUT(n24969), .C0(n1731), .Z(n14662));
    LUT4 i2_4_lut_adj_247 (.A(n26540), .B(n28548), .C(register_addr[0]), 
         .D(prev_select), .Z(n8273)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_247.init = 16'h0008;
    LUT4 i5422_3_lut (.A(debug_c_7), .B(n1278[3]), .C(n1278[2]), .Z(n11426)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5422_3_lut.init = 16'h5454;
    LUT4 i2_4_lut_adj_248 (.A(n28474), .B(n28477), .C(n26399), .D(prev_select_adj_177), 
         .Z(n3452)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_4_lut_adj_248.init = 16'h0020;
    LUT4 i2_4_lut_adj_249 (.A(databus[4]), .B(n5_adj_377), .C(n1278[13]), 
         .D(n26365), .Z(n24660)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_249.init = 16'hffec;
    LUT4 select_1894_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1278[4]), 
         .C(rx_data[4]), .D(n26579), .Z(n5_adj_377)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_250 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [1]), 
         .Z(n26384)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_250.init = 16'h2020;
    LUT4 i13320_3_lut_4_lut (.A(n28455), .B(n1278[14]), .C(n9_adj_353), 
         .D(sendcount[0]), .Z(n18[0])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i13320_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i2_4_lut_adj_251 (.A(databus[3]), .B(n5_adj_378), .C(n1278[13]), 
         .D(n26364), .Z(n24661)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_251.init = 16'hffec;
    LUT4 i2_2_lut (.A(n1278[17]), .B(n1278[9]), .Z(n8_c)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1278[4]), .B(n28580), .C(bufcount[0]), 
         .D(n28447), .Z(n24846)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hd222;
    LUT4 i1_4_lut_adj_252 (.A(n28534), .B(n1278[18]), .C(n8_adj_379), 
         .D(n1278[6]), .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_252.init = 16'hfffe;
    LUT4 select_1894_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1278[4]), 
         .C(rx_data[3]), .D(n26579), .Z(n5_adj_378)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n28574), .B(n28511), .C(n4_adj_311), 
         .D(n28585), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i916_3_lut (.A(n1278[5]), .B(n28485), .C(n1278[10]), .Z(n2592)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i916_3_lut.init = 16'hc8c8;
    LUT4 i2_4_lut_adj_253 (.A(databus[2]), .B(n5_adj_380), .C(n1278[13]), 
         .D(n26362), .Z(n24659)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_253.init = 16'hffec;
    LUT4 select_1894_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1278[4]), 
         .C(rx_data[2]), .D(n26579), .Z(n5_adj_380)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_254 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n26578)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_254.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_4_lut_adj_255 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][14] ), .D(n28542), .Z(n26079)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_255.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_256 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][12] ), .D(n28542), .Z(n26098)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_256.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_257 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n26579)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_257.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_258 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][10] ), .D(n28542), .Z(n26081)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_258.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_259 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][7] ), .D(n28542), .Z(n26090)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_259.init = 16'h1000;
    LUT4 i2_4_lut_adj_260 (.A(databus[1]), .B(n5_adj_381), .C(n1278[13]), 
         .D(n26361), .Z(n24662)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_260.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_261 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][11] ), .D(n28542), .Z(n26083)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_261.init = 16'h1000;
    LUT4 i20_2_lut_rep_327_3_lut_4_lut (.A(select[4]), .B(n28565), .C(rw), 
         .D(n28519), .Z(n28448)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i20_2_lut_rep_327_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_331_3_lut_4_lut (.A(select[4]), .B(n28565), .C(n28578), 
         .D(register_addr_c[5]), .Z(n28452)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_331_3_lut_4_lut.init = 16'h0008;
    LUT4 equal_182_i4_2_lut_rep_456 (.A(bufcount[1]), .B(bufcount[2]), .Z(n28577)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam equal_182_i4_2_lut_rep_456.init = 16'heeee;
    LUT4 i2612_2_lut_rep_375_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n28496)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i2612_2_lut_rep_375_3_lut.init = 16'hfefe;
    LUT4 select_1894_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1278[4]), 
         .C(rx_data[1]), .D(n26579), .Z(n5_adj_381)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_262 (.A(n1278[3]), .B(n28486), .C(\buffer[5] [0]), 
         .Z(n26383)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_262.init = 16'h2020;
    LUT4 i1_2_lut_adj_263 (.A(register_addr[0]), .B(\control_reg[7] ), .Z(n7685)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_263.init = 16'h4444;
    LUT4 i2_3_lut_rep_457 (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr_c[3]), .Z(n28578)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_457.init = 16'hfefe;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n28574), .B(n28511), .C(n4_adj_302), 
         .D(n28588), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i259_2_lut_rep_393_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr_c[3]), .D(register_addr_c[5]), .Z(n28514)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i259_2_lut_rep_393_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_264 (.A(register_addr[0]), .B(\control_reg[7]_adj_181 ), 
         .Z(n7694)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_264.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_265 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][6] ), .D(n28542), .Z(n26088)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_265.init = 16'h1000;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n28574), .B(n28511), .C(n4_adj_301), 
         .D(n28597), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_adj_266 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [7]), 
         .Z(n26382)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_266.init = 16'h2020;
    LUT4 i1_2_lut_4_lut_adj_267 (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr_c[3]), .D(prev_select), .Z(n151)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_267.init = 16'hfffe;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n28574), .B(n28511), .C(n4_adj_300), 
         .D(n28603), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i2_4_lut_adj_268 (.A(databus[0]), .B(n5_adj_383), .C(n1278[13]), 
         .D(n26388), .Z(n24808)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_268.init = 16'hffec;
    LUT4 select_1894_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1278[4]), 
         .C(rx_data[0]), .D(n26579), .Z(n5_adj_383)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_398_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr_c[3]), .D(register_addr_c[5]), .Z(n28519)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_398_4_lut.init = 16'h0100;
    LUT4 n27980_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n28567), .C(n28615), 
         .D(n27980), .Z(n27981)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n27980_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 i885_2_lut_rep_458 (.A(escape), .B(debug_c_7), .Z(n28579)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i885_2_lut_rep_458.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_269 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][5] ), .D(n28542), .Z(n26096)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_269.init = 16'h1000;
    PFUMX i20876 (.BLUT(n28583), .ALUT(n28584), .C0(sendcount[0]), .Z(n28585));
    LUT4 i1_2_lut_3_lut_adj_270 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [6]), 
         .Z(n26381)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_270.init = 16'h2020;
    LUT4 i1_4_lut_adj_271 (.A(n1278[4]), .B(\buffer[1] [7]), .C(n11_adj_384), 
         .D(n14_c), .Z(n25655)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_271.init = 16'heca0;
    LUT4 i1_4_lut_adj_272 (.A(n1278[4]), .B(\buffer[1] [6]), .C(n11_adj_385), 
         .D(n14_c), .Z(n25679)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_272.init = 16'heca0;
    LUT4 i2_3_lut_rep_326_4_lut (.A(escape), .B(debug_c_7), .C(n28486), 
         .D(n1278[4]), .Z(n28447)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_326_4_lut.init = 16'hffbf;
    LUT4 i1_2_lut_3_lut_4_lut_adj_273 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][9] ), .D(n28542), .Z(n26077)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_273.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_274 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [5]), 
         .Z(n26380)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_274.init = 16'h2020;
    LUT4 i1_3_lut_rep_459 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n28580)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_rep_459.init = 16'hecec;
    LUT4 i2_2_lut_rep_388_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1278[4]), .Z(n28509)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_388_4_lut.init = 16'hecff;
    LUT4 i1_4_lut_adj_275 (.A(n1278[4]), .B(\buffer[1] [5]), .C(n11_adj_386), 
         .D(n14_c), .Z(n25677)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_275.init = 16'heca0;
    LUT4 i1_4_lut_adj_276 (.A(n1278[4]), .B(\buffer[1] [4]), .C(n11_adj_387), 
         .D(n14_c), .Z(n25657)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_276.init = 16'heca0;
    LUT4 i1_2_lut_4_lut_adj_277 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1278[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_277.init = 16'hec00;
    LUT4 i1_2_lut_3_lut_4_lut_adj_278 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][8] ), .D(n28542), .Z(n26076)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_278.init = 16'h1000;
    LUT4 i1_4_lut_adj_279 (.A(n1278[4]), .B(\buffer[1] [3]), .C(n11_adj_388), 
         .D(n14_c), .Z(n25741)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_279.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_adj_280 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [4]), 
         .Z(n26379)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_280.init = 16'h2020;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n28577), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_384)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_281 (.A(bufcount[0]), .B(n28577), .C(\buffer[1] [6]), 
         .D(rx_data[6]), .Z(n11_adj_385)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_281.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_282 (.A(bufcount[0]), .B(n28577), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_386)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_282.init = 16'hf2d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_283 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][13] ), .D(n28542), .Z(n26085)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_283.init = 16'h1000;
    LUT4 i1_4_lut_adj_284 (.A(n1278[4]), .B(\buffer[1] [2]), .C(n11_adj_389), 
         .D(n14_c), .Z(n25729)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_284.init = 16'heca0;
    LUT4 i1_4_lut_adj_285 (.A(n1278[4]), .B(debug_c_7), .C(n1278[2]), 
         .D(n26299), .Z(n25771)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_285.init = 16'heeea;
    LUT4 i24_3_lut_4_lut_adj_286 (.A(bufcount[0]), .B(n28577), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_387)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_286.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_287 (.A(bufcount[0]), .B(n28577), .C(rx_data[3]), 
         .D(\buffer[1] [3]), .Z(n11_adj_388)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_287.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_adj_288 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [3]), 
         .Z(n26372)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_288.init = 16'h2020;
    LUT4 i24_3_lut_4_lut_adj_289 (.A(bufcount[0]), .B(n28577), .C(rx_data[2]), 
         .D(\buffer[1] [2]), .Z(n11_adj_389)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_289.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_290 (.A(bufcount[0]), .B(n28577), .C(rx_data[1]), 
         .D(\buffer[1] [1]), .Z(n11_adj_390)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_290.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_291 (.A(bufcount[0]), .B(n28577), .C(\buffer[1] [0]), 
         .D(rx_data[0]), .Z(n11_adj_391)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_291.init = 16'hf2d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_292 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][4] ), .D(n28542), .Z(n26100)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_292.init = 16'h1000;
    LUT4 i1_2_lut_rep_338_3_lut (.A(register_addr_c[5]), .B(n28578), .C(register_addr_c[4]), 
         .Z(n28459)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_338_3_lut.init = 16'hfefe;
    LUT4 n28486_bdd_4_lut (.A(bufcount[1]), .B(n1278[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n29190)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n28486_bdd_4_lut.init = 16'h0080;
    LUT4 i1_4_lut_adj_293 (.A(n1278[4]), .B(\buffer[1] [1]), .C(n11_adj_390), 
         .D(n14_c), .Z(n25743)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_293.init = 16'heca0;
    LUT4 n28486_bdd_4_lut_21199 (.A(n28486), .B(n28579), .C(n1278[0]), 
         .D(n1278[3]), .Z(n29188)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C)) */ ;
    defparam n28486_bdd_4_lut_21199.init = 16'hdd0f;
    LUT4 i1_2_lut_rep_310_3_lut_4_lut (.A(register_addr_c[5]), .B(n28578), 
         .C(register_addr[2]), .D(register_addr_c[4]), .Z(n28431)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_310_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_319_3_lut_4_lut (.A(register_addr_c[5]), .B(n28578), 
         .C(register_addr[1]), .D(register_addr_c[4]), .Z(n28440)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_319_3_lut_4_lut.init = 16'hfffe;
    LUT4 i8793_3_lut_4_lut (.A(register_addr[2]), .B(n28459), .C(n11), 
         .D(n12585), .Z(n14798)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i8793_3_lut_4_lut.init = 16'hef00;
    LUT4 i1_4_lut_adj_294 (.A(n1278[4]), .B(\buffer[1] [0]), .C(n11_adj_391), 
         .D(n14_c), .Z(n25693)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_294.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_295 (.A(register_addr_c[5]), .B(n28578), 
         .C(register_addr[1]), .D(n28565), .Z(n26514)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_295.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_296 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][15] ), .D(n28542), .Z(n26087)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_296.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_297 (.A(register_addr_c[5]), .B(n28578), 
         .C(register_addr[1]), .D(n28565), .Z(n26540)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_297.init = 16'h1000;
    LUT4 i1_2_lut_adj_298 (.A(register_addr[0]), .B(\control_reg[7]_adj_182 ), 
         .Z(n7703)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_298.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_299 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [2]), 
         .Z(n26378)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_299.init = 16'h2020;
    LUT4 i20_2_lut_rep_330_3_lut_4_lut (.A(register_addr_c[5]), .B(n28578), 
         .C(n30468), .D(n28517), .Z(n28451)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i20_2_lut_rep_330_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_300 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [1]), 
         .Z(n26377)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_300.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_301 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][16] ), .D(n28542), .Z(n26084)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_301.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_302 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][17] ), .D(n28542), .Z(n26094)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_302.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_303 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][18] ), .D(n28542), .Z(n26095)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_303.init = 16'h1000;
    LUT4 i1_4_lut_adj_304 (.A(n1278[4]), .B(\buffer[0] [7]), .C(n11_adj_393), 
         .D(n14_c), .Z(n25695)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_304.init = 16'heca0;
    LUT4 i1_2_lut_adj_305 (.A(register_addr[1]), .B(\steps_reg[5] ), .Z(n14)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_305.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_306 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][19] ), .D(n28542), .Z(n26093)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_306.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_307 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][20] ), .D(n28542), .Z(n26091)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_307.init = 16'h1000;
    FD1S3IX state_FSM_i21 (.D(n11252), .CK(debug_c_c), .CD(n30473), .Q(n1278[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_308 (.A(n15_c), .B(n1278[3]), .C(n1278[0]), .D(n26738), 
         .Z(n26299)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_308.init = 16'h50dc;
    LUT4 i1_4_lut_adj_309 (.A(n1278[4]), .B(\buffer[0] [6]), .C(n11_adj_395), 
         .D(n14_c), .Z(n25651)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_309.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_310 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][21] ), .D(n28542), .Z(n26092)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_310.init = 16'h1000;
    LUT4 Select_3927_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[21]_adj_183 ), 
         .D(rw), .Z(n1_adj_184)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3927_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_359_3_lut_4_lut (.A(n28547), .B(select[4]), .C(n28578), 
         .D(register_addr_c[5]), .Z(n28480)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_359_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_311 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][22] ), .D(n28542), .Z(n26080)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_311.init = 16'h1000;
    LUT4 n26402_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n27600)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n26402_bdd_4_lut.init = 16'h4001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_312 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][23] ), .D(n28542), .Z(n26086)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_312.init = 16'h1000;
    LUT4 i20_2_lut_rep_337_3_lut_4_lut (.A(n28547), .B(select[4]), .C(rw), 
         .D(n28519), .Z(n28458)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i20_2_lut_rep_337_3_lut_4_lut.init = 16'h4000;
    FD1S3IX state_FSM_i20 (.D(n10029), .CK(debug_c_c), .CD(n30473), .Q(n1278[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n25785), .CK(debug_c_c), .CD(n30473), .Q(n1278[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n11254), .CK(debug_c_c), .CD(n30473), .Q(n1278[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n10023), .CK(debug_c_c), .CD(n30473), .Q(n1278[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1390), .CK(debug_c_c), .CD(n30473), .Q(n1278[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1389), .CK(debug_c_c), .CD(n30473), .Q(n1278[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1278[12]), .CK(debug_c_c), .CD(n30473), 
            .Q(n1278[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1278[11]), .CK(debug_c_c), .CD(n30473), 
            .Q(n1278[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1278[10]), .CK(debug_c_c), .CD(n30473), 
            .Q(n1278[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1383), .CK(debug_c_c), .CD(n30473), .Q(n1278[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1278[8]), .CK(debug_c_c), .CD(n30473), 
            .Q(n1278[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1278[7]), .CK(debug_c_c), .CD(n30473), .Q(n1278[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    LUT4 mux_1703_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n5020), 
         .Z(n5011[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1703_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_313 (.A(n1278[4]), .B(\buffer[0] [5]), .C(n11_adj_398), 
         .D(n14_c), .Z(n25727)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_313.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_adj_314 (.A(n1278[3]), .B(n28486), .C(\buffer[4] [0]), 
         .Z(n26376)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_314.init = 16'h2020;
    FD1S3IX state_FSM_i8 (.D(n1278[6]), .CK(debug_c_c), .CD(n30473), .Q(n1278[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1278[5]), .CK(debug_c_c), .CD(n30473), .Q(n1278[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n26464), .CK(debug_c_c), .CD(n30473), .Q(n1278[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n26298), .CK(debug_c_c), .CD(n30473), .Q(n1278[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n11426), .CK(debug_c_c), .CD(n30473), .Q(n1278[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n25771), .CK(debug_c_c), .CD(n30473), .Q(n1278[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i2 (.D(n25885), .CK(debug_c_c), .CD(n30473), .Q(n1278[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    LUT4 i24_3_lut_4_lut_adj_315 (.A(bufcount[0]), .B(n28577), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_adj_306)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_315.init = 16'hf1e0;
    LUT4 i20044_3_lut (.A(n12121), .B(escape), .C(n15_c), .Z(n26738)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i20044_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_316 (.A(n1278[4]), .B(\buffer[0] [4]), .C(n11_adj_399), 
         .D(n14_c), .Z(n25659)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_316.init = 16'heca0;
    LUT4 i24_3_lut_4_lut_adj_317 (.A(bufcount[0]), .B(n28577), .C(rx_data[7]), 
         .D(\buffer[0] [7]), .Z(n11_adj_393)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_317.init = 16'hfe10;
    LUT4 i1_2_lut_3_lut_4_lut_adj_318 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][24] ), .D(n28542), .Z(n26078)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_318.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_319 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][25] ), .D(n28542), .Z(n26082)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_319.init = 16'h1000;
    LUT4 i24_3_lut_4_lut_adj_320 (.A(bufcount[0]), .B(n28577), .C(\buffer[0] [6]), 
         .D(rx_data[6]), .Z(n11_adj_395)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_320.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_321 (.A(n1278[4]), .B(\buffer[0] [3]), .C(n11_adj_400), 
         .D(n14_c), .Z(n25681)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_321.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_322 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][26] ), .D(n28542), .Z(n26089)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_322.init = 16'h1000;
    LUT4 i24_3_lut_4_lut_adj_323 (.A(bufcount[0]), .B(n28577), .C(rx_data[5]), 
         .D(\buffer[0] [5]), .Z(n11_adj_398)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_323.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_324 (.A(bufcount[0]), .B(n28577), .C(\buffer[0] [4]), 
         .D(rx_data[4]), .Z(n11_adj_399)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_324.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_325 (.A(n1278[4]), .B(\buffer[0] [2]), .C(n11_adj_401), 
         .D(n14_c), .Z(n25675)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_325.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_326 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][27] ), .D(n28542), .Z(n26102)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_326.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_327 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][28] ), .D(n28542), .Z(n26097)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_327.init = 16'h1000;
    LUT4 i24_3_lut_4_lut_adj_328 (.A(bufcount[0]), .B(n28577), .C(rx_data[3]), 
         .D(\buffer[0] [3]), .Z(n11_adj_400)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_328.init = 16'hfe10;
    LUT4 i1_2_lut_3_lut_adj_329 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [7]), 
         .Z(n26375)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_329.init = 16'h2020;
    LUT4 i24_3_lut_4_lut_adj_330 (.A(bufcount[0]), .B(n28577), .C(\buffer[0] [2]), 
         .D(rx_data[2]), .Z(n11_adj_401)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_330.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_331 (.A(bufcount[0]), .B(n28577), .C(\buffer[0] [1]), 
         .D(rx_data[1]), .Z(n11_adj_402)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_331.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_332 (.A(n1278[4]), .B(\buffer[0] [1]), .C(n11_adj_402), 
         .D(n14_c), .Z(n25673)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_332.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_333 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][29] ), .D(n28542), .Z(n26099)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_333.init = 16'h1000;
    LUT4 i8292_4_lut (.A(escape), .B(n12121), .C(n6_adj_403), .D(n1278[3]), 
         .Z(n9903)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i8292_4_lut.init = 16'h1aaa;
    LUT4 i1_2_lut_3_lut_4_lut_adj_334 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][30] ), .D(n28542), .Z(n26103)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_334.init = 16'h1000;
    LUT4 i2_2_lut_adj_335 (.A(debug_c_7), .B(n28485), .Z(n6_adj_403)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_335.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_336 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [6]), 
         .Z(n26371)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_336.init = 16'h2020;
    LUT4 i3_4_lut_adj_337 (.A(n1278[7]), .B(n1278[2]), .C(n28535), .D(n1278[10]), 
         .Z(n8_adj_379)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_337.init = 16'hfffe;
    LUT4 i2_4_lut_adj_338 (.A(n28419), .B(n28477), .C(n183), .D(prev_select_adj_176), 
         .Z(n3626)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_338.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_339 (.A(register_addr_c[5]), .B(n28578), 
         .C(register_addr[1]), .D(n28547), .Z(n26489)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_339.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_adj_340 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [5]), 
         .Z(n26373)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_340.init = 16'h2020;
    LUT4 i1_2_lut_rep_355_3_lut_4_lut (.A(register_addr_c[5]), .B(n28578), 
         .C(n28565), .D(select[4]), .Z(n28476)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_355_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_366_3_lut_4_lut (.A(register_addr_c[5]), .B(n28578), 
         .C(select[4]), .D(n28547), .Z(n28487)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_366_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_341 (.A(register_addr_c[5]), .B(n28578), 
         .C(register_addr[1]), .D(n28565), .Z(n26437)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_341.init = 16'h0200;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_368)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_4_lut_adj_342 (.A(register_addr_c[5]), .B(n28578), 
         .C(register_addr[1]), .D(n28565), .Z(n26439)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_342.init = 16'h2000;
    LUT4 i1_4_lut_adj_343 (.A(n28496), .B(debug_c_7), .C(n12374), .D(n8_adj_404), 
         .Z(n25885)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_343.init = 16'hdc50;
    LUT4 i1_2_lut_3_lut_4_lut_adj_344 (.A(register_addr_c[5]), .B(n28578), 
         .C(n28547), .D(register_addr[1]), .Z(n233)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_344.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_345 (.A(register_addr[2]), .B(n28459), 
         .C(\register[2][31] ), .D(n28542), .Z(n26101)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_345.init = 16'h1000;
    LUT4 i2_4_lut_adj_346 (.A(n28578), .B(n28565), .C(prev_select_adj_185), 
         .D(n28497), .Z(n26396)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i2_4_lut_adj_346.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_347 (.A(register_addr[2]), .B(n28459), 
         .C(n183), .D(n12585), .Z(n8472)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_347.init = 16'h1000;
    LUT4 i1_2_lut_adj_348 (.A(register_addr[1]), .B(\steps_reg[6] ), .Z(n13)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_348.init = 16'h8888;
    LUT4 i1_3_lut (.A(n15_c), .B(n1278[1]), .C(n1278[0]), .Z(n8_adj_404)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_adj_349 (.A(register_addr[1]), .B(\steps_reg[3] ), .Z(n12)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_349.init = 16'h8888;
    LUT4 i1_2_lut_adj_350 (.A(register_addr[1]), .B(register_addr[0]), .Z(n183)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_350.init = 16'h8888;
    LUT4 Select_3929_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[20]_adj_186 ), 
         .D(rw), .Z(n1_adj_187)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3929_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_351 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [4]), 
         .Z(n26374)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_351.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_352 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [3]), 
         .Z(n26370)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_352.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_353 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [2]), 
         .Z(n26369)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_353.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_354 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [1]), 
         .Z(n26368)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_354.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_355 (.A(n1278[3]), .B(n28486), .C(\buffer[3] [0]), 
         .Z(n26359)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_355.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_356 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [7]), 
         .Z(n26358)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_356.init = 16'h2020;
    LUT4 i4_4_lut_adj_357 (.A(n1278[4]), .B(n26631), .C(n1278[20]), .D(n6), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_357.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_358 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [6]), 
         .Z(n26367)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_358.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_359 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [5]), 
         .Z(n26366)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_359.init = 16'h2020;
    LUT4 i13150_2_lut (.A(bufcount[0]), .B(n1278[0]), .Z(n14663)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i13150_2_lut.init = 16'h2222;
    LUT4 Select_3931_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[19]_adj_188 ), 
         .D(n30468), .Z(n1_adj_189)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3931_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_360 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [4]), 
         .Z(n26365)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_360.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_361 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [3]), 
         .Z(n26364)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_361.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_362 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [2]), 
         .Z(n26362)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_362.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_363 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [1]), 
         .Z(n26361)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_363.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_364 (.A(n1278[3]), .B(n28486), .C(\buffer[2] [0]), 
         .Z(n26388)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_364.init = 16'h2020;
    LUT4 i20328_2_lut_2_lut (.A(n28485), .B(n8417), .Z(n13149)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i20328_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_1703_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n5020), 
         .Z(n5011[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1703_i3_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_365 (.A(n1278[16]), .B(n1278[19]), .Z(n2029)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_365.init = 16'heeee;
    LUT4 Select_3933_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[18]_adj_190 ), 
         .D(rw), .Z(n1_adj_191)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3933_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3935_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[17]_adj_192 ), 
         .D(rw), .Z(n1_adj_193)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3935_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_366 (.A(n28466), .B(n28542), .C(n28547), .D(n28477), 
         .Z(n12981)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i1_2_lut_4_lut_adj_366.init = 16'hff08;
    LUT4 Select_3937_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[16]_adj_194 ), 
         .D(n30468), .Z(n1_adj_195)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3937_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_367 (.A(register_addr[1]), .B(n28459), 
         .C(register_addr[2]), .D(register_addr[0]), .Z(n15)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_367.init = 16'hffef;
    LUT4 i13024_2_lut_3_lut_4_lut (.A(register_addr_c[4]), .B(n28514), .C(register_addr[1]), 
         .D(register_addr[2]), .Z(n8336)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i13024_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_368 (.A(register_addr_c[4]), .B(n28514), 
         .C(register_addr[0]), .D(register_addr[2]), .Z(n4_adj_196)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_368.init = 16'hfffe;
    LUT4 i2_4_lut_adj_369 (.A(n26454), .B(n28468), .C(n28578), .D(prev_select_adj_176), 
         .Z(n12580)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_369.init = 16'h0002;
    LUT4 i20361_2_lut_3_lut_3_lut_4_lut_4_lut (.A(register_addr[1]), .B(n28459), 
         .C(register_addr[0]), .D(register_addr[2]), .Z(n62)) /* synthesis lut_function=(!(A (B+(D))+!A (B+(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i20361_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h0133;
    LUT4 i1_2_lut_3_lut_4_lut_adj_370 (.A(register_addr[1]), .B(n28459), 
         .C(register_addr[2]), .D(register_addr[0]), .Z(n15_adj_197)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_370.init = 16'hfffe;
    LUT4 n27504_bdd_2_lut_3_lut_4_lut (.A(register_addr_c[4]), .B(n28514), 
         .C(n27504), .D(register_addr[2]), .Z(n27505)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n27504_bdd_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 n27502_bdd_2_lut_3_lut_4_lut (.A(register_addr_c[4]), .B(n28514), 
         .C(n27502), .D(register_addr[2]), .Z(n27503)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n27502_bdd_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_298_3_lut_4_lut (.A(register_addr_c[4]), .B(n28514), 
         .C(n28548), .D(register_addr[2]), .Z(n28419)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_298_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_371 (.A(n1278[6]), .B(n1278[11]), .Z(n1731)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_371.init = 16'heeee;
    LUT4 i3_4_lut_adj_372 (.A(\buffer[0] [3]), .B(\buffer[0] [5]), .C(\buffer[0] [4]), 
         .D(\buffer[0] [6]), .Z(n12_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i3_4_lut_adj_372.init = 16'hfffe;
    LUT4 i20336_2_lut_rep_304_3_lut_4_lut (.A(register_addr_c[4]), .B(n28514), 
         .C(register_addr[1]), .D(register_addr[2]), .Z(n28425)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i20336_2_lut_rep_304_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_3_lut_rep_318_4_lut (.A(register_addr_c[4]), .B(n28514), .C(n183), 
         .D(register_addr[2]), .Z(n28439)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_3_lut_rep_318_4_lut.init = 16'hfeee;
    LUT4 i20371_4_lut (.A(\buffer[0] [2]), .B(n12_c), .C(\buffer[0] [0]), 
         .D(\buffer[0] [1]), .Z(n24909)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i20371_4_lut.init = 16'h2000;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_367)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i43_1_lut_3_lut_4_lut (.A(register_addr_c[4]), .B(n28514), .C(n183), 
         .D(register_addr[2]), .Z(n176)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i43_1_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 Select_3939_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[15]_adj_198 ), 
         .D(n30468), .Z(n1_adj_199)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3939_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i20331_4_lut (.A(\buffer[0] [2]), .B(\buffer[0] [1]), .C(\buffer[0] [0]), 
         .D(n12_c), .Z(n24969)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i20331_4_lut.init = 16'h0004;
    LUT4 i4_4_lut_adj_373 (.A(n1278[10]), .B(n8_adj_423), .C(n1278[13]), 
         .D(n26631), .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_373.init = 16'hfffe;
    LUT4 i3_3_lut (.A(n1278[9]), .B(n1278[11]), .C(n1278[8]), .Z(n8_adj_423)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_3_lut.init = 16'hfefe;
    LUT4 Select_3941_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[14]_adj_200 ), 
         .D(n30468), .Z(n1_adj_201)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3941_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1703_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n5020), 
         .Z(n5011[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1703_i2_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_adj_365)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 Select_3945_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[12]_adj_202 ), 
         .D(n30468), .Z(n1_adj_203)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3945_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3953_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[8]_adj_204 ), 
         .D(n30468), .Z(n1_adj_205)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3953_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_374 (.A(n28419), .B(prev_select_adj_176), .C(n28542), 
         .D(n28477), .Z(n12647)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_374.init = 16'hff20;
    LUT4 rx_data_2__bdd_4_lut_21148 (.A(rx_data[2]), .B(rx_data[3]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n27797)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_2__bdd_4_lut_21148.init = 16'h6001;
    LUT4 i13164_4_lut (.A(sendcount[3]), .B(n9_adj_353), .C(sendcount[2]), 
         .D(n28566), .Z(n19[3])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(271[10:37])
    defparam i13164_4_lut.init = 16'h4888;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n28449), .CD(n14807), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n28449), .CD(n14807), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n28449), .CD(n14807), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n28449), .CD(n14807), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n12642), .CD(n14803), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    LUT4 mux_500_i5_3_lut (.A(n2537), .B(esc_data[4]), .C(n1278[18]), 
         .Z(n2020[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_500_i5_3_lut.init = 16'hcaca;
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n12642), .CD(n14803), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n12642), .CD(n14803), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n12642), .CD(n14803), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 mux_500_i4_3_lut (.A(n2537), .B(esc_data[3]), .C(n1278[18]), 
         .Z(n2020[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_500_i4_3_lut.init = 16'hcaca;
    LUT4 mux_500_i2_3_lut (.A(n2537), .B(esc_data[1]), .C(n1278[18]), 
         .Z(n2020[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_500_i2_3_lut.init = 16'hcaca;
    LUT4 sendcount_1__bdd_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(sendcount[3]), 
         .D(sendcount[2]), .Z(n27814)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_1__bdd_4_lut.init = 16'h6aaa;
    LUT4 Select_3949_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[10]_adj_206 ), 
         .D(rw), .Z(n1_adj_207)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3949_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3909_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[30]_adj_208 ), 
         .D(n30468), .Z(n1_adj_209)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3909_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_375 (.A(databus[31]), .B(n5_adj_434), .C(n1278[13]), 
         .D(n26363), .Z(n24764)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_375.init = 16'hffec;
    LUT4 select_1894_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1278[4]), 
         .C(rx_data[7]), .D(n26570), .Z(n5_adj_434)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1894_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 sendcount_4__bdd_3_lut (.A(sendcount[4]), .B(n27814), .C(\sendcount[1] ), 
         .Z(n27815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_376 (.A(n28519), .B(n28510), .C(prev_select_adj_185), 
         .D(n28477), .Z(n12599)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_376.init = 16'h0008;
    LUT4 Select_3951_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[9]_adj_210 ), 
         .D(rw), .Z(n1_adj_211)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3951_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX rw_498_rep_463 (.D(n1278[10]), .SP(n2592), .CK(debug_c_c), 
            .Q(n30468));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_463.GSR = "ENABLED";
    LUT4 Select_3947_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[11]_adj_212 ), 
         .D(rw), .Z(n1_adj_213)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3947_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3943_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[13]_adj_214 ), 
         .D(rw), .Z(n1_adj_215)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3943_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_324_4_lut (.A(n28497), .B(n28578), .C(prev_select_adj_177), 
         .D(n28468), .Z(n28445)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i1_2_lut_rep_324_4_lut.init = 16'h0002;
    LUT4 Select_3915_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[27]_adj_216 ), 
         .D(n30468), .Z(n1_adj_217)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3915_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3913_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[28]_adj_218 ), 
         .D(n30468), .Z(n1_adj_219)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3913_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3907_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[31]_adj_220 ), 
         .D(n30468), .Z(n1_adj_221)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3907_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3911_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[29]_adj_222 ), 
         .D(rw), .Z(n1_adj_223)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3911_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3960_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[1] ), 
         .D(rw), .Z(n1_adj_224)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3960_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3917_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[26]_adj_225 ), 
         .D(n30468), .Z(n1_adj_226)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3917_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_377 (.A(register_addr[0]), .B(n28500), 
         .C(n28477), .D(n28466), .Z(n12995)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_377.init = 16'hf1f0;
    PFUMX i20721 (.BLUT(n27981), .ALUT(n27976), .C0(n5020), .Z(n27982));
    LUT4 i5250_3_lut (.A(busy), .B(n1278[20]), .C(n1278[19]), .Z(n11252)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5250_3_lut.init = 16'ha8a8;
    LUT4 i4030_3_lut (.A(n1278[19]), .B(n1278[18]), .C(busy), .Z(n10029)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4030_3_lut.init = 16'hcece;
    LUT4 i2_4_lut_adj_378 (.A(n38), .B(busy), .C(n27601), .D(n1278[17]), 
         .Z(n25785)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_378.init = 16'hfbfa;
    LUT4 i1_4_lut_adj_379 (.A(n1278[15]), .B(esc_data[7]), .C(n8_adj_452), 
         .D(esc_data[0]), .Z(n38)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_379.init = 16'ha8aa;
    LUT4 Select_3919_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[25]_adj_227 ), 
         .D(n30468), .Z(n1_adj_228)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3919_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3921_i1_2_lut_3_lut_4_lut (.A(n28519), .B(n28510), .C(\read_value[24]_adj_229 ), 
         .D(n30468), .Z(n1_adj_230)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3921_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_380 (.A(n35), .B(esc_data[5]), .C(n55), .D(esc_data[6]), 
         .Z(n8_adj_452)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_380.init = 16'hfffe;
    LUT4 i1_4_lut_adj_381 (.A(esc_data[4]), .B(esc_data[3]), .C(esc_data[1]), 
         .D(esc_data[2]), .Z(n35)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_381.init = 16'h5f4c;
    LUT4 i51_4_lut (.A(esc_data[2]), .B(esc_data[3]), .C(esc_data[4]), 
         .D(esc_data[1]), .Z(n55)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i51_4_lut.init = 16'h9998;
    LUT4 i5251_3_lut (.A(busy), .B(n1278[17]), .C(n1278[16]), .Z(n11254)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5251_3_lut.init = 16'ha8a8;
    LUT4 i4024_3_lut (.A(n1278[16]), .B(n2537), .C(busy), .Z(n10023)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4024_3_lut.init = 16'hcece;
    LUT4 i449_2_lut (.A(n5020), .B(n1278[14]), .Z(n1390)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i449_2_lut.init = 16'h4444;
    LUT4 reduce_or_447_i1_3_lut (.A(busy), .B(n1278[13]), .C(n1278[20]), 
         .Z(n1389)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_447_i1_3_lut.init = 16'hdcdc;
    LUT4 i1_2_lut_adj_382 (.A(register_addr[1]), .B(\steps_reg[7] ), .Z(n12_adj_231)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_382.init = 16'h8888;
    LUT4 i4_4_lut_adj_383 (.A(rx_data[2]), .B(n26319), .C(rx_data[5]), 
         .D(n6_adj_458), .Z(n12374)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i4_4_lut_adj_383.init = 16'h0800;
    LUT4 i2_4_lut_adj_384 (.A(escape), .B(n12174), .C(debug_c_7), .D(n28581), 
         .Z(n26319)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2_4_lut_adj_384.init = 16'h0040;
    LUT4 i1_2_lut_adj_385 (.A(n1278[3]), .B(rx_data[0]), .Z(n6_adj_458)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_adj_385.init = 16'h8888;
    PFUMX i20896 (.BLUT(n28613), .ALUT(n28614), .C0(sendcount[0]), .Z(n28615));
    PFUMX i20894 (.BLUT(n28610), .ALUT(n28611), .C0(sendcount[3]), .Z(n5020));
    PFUMX i20892 (.BLUT(n28607), .ALUT(n28608), .C0(sendcount[0]), .Z(n28609));
    PFUMX i20890 (.BLUT(n28604), .ALUT(n28605), .C0(sendcount[0]), .Z(n28606));
    PFUMX i20888 (.BLUT(n28601), .ALUT(n28602), .C0(sendcount[0]), .Z(n28603));
    PFUMX i20886 (.BLUT(n28598), .ALUT(n28599), .C0(sendcount[0]), .Z(n28600));
    PFUMX i20884 (.BLUT(n28595), .ALUT(n28596), .C0(sendcount[0]), .Z(n28597));
    PFUMX i20882 (.BLUT(n28592), .ALUT(n28593), .C0(n28447), .Z(n28594));
    PFUMX i20878 (.BLUT(n28586), .ALUT(n28587), .C0(sendcount[0]), .Z(n28588));
    \UARTTransmitter(baud_div=12)  uart_output (.n30473(n30473), .tx_data({tx_data}), 
            .send(send), .\reset_count[7] (\reset_count[7] ), .\reset_count[6] (\reset_count[6] ), 
            .\reset_count[5] (\reset_count[5] ), .n24551(n24551), .n28485(n28485), 
            .n4(n4_c), .n5020(n5020), .n1296(n1278[14]), .n12642(n12642), 
            .n1293(n1278[17]), .n1290(n1278[20]), .n24779(n24779), .n9969(n9969), 
            .busy(busy), .GND_net(GND_net), .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_c(debug_c_c), .n28485(n28485), 
            .rx_data({rx_data}), .n30473(n30473), .n28457(n28457), .debug_c_7(debug_c_7), 
            .n9970_c(n9970_c), .n28581(n28581), .n28518(n28518), .n28486(n28486), 
            .n15(n15_c), .n12121(n12121), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (n30473, tx_data, send, \reset_count[7] , 
            \reset_count[6] , \reset_count[5] , n24551, n28485, n4, 
            n5020, n1296, n12642, n1293, n1290, n24779, n9969, 
            busy, GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input n30473;
    input [7:0]tx_data;
    input send;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n24551;
    input n28485;
    input n4;
    input n5020;
    input n1296;
    output n12642;
    input n1293;
    input n1290;
    output n24779;
    output n9969;
    output busy;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27868, n27867;
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n27869;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n8399, n12687, n26334, n26829, n26830, n26831, n17, n17_adj_299, 
        n28553, n11, n25937, n25763, n7, n10, n104, n10070, 
        n13549, n19307, n26766, n2;
    
    PFUMX i20683 (.BLUT(n27868), .ALUT(n27867), .C0(state[2]), .Z(n27869));
    FD1S3IX state__i0 (.D(n27869), .CK(bclk), .CD(n30473), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n8399), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n8399), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n8399), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n8399), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n8399), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n8399), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n8399), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n8399), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n26334), .SP(n12687), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    PFUMX i20135 (.BLUT(n26829), .ALUT(n26830), .C0(state[1]), .Z(n26831));
    LUT4 state_2__bdd_2_lut (.A(state[0]), .B(state[3]), .Z(n27867)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_2__bdd_2_lut.init = 16'h1111;
    LUT4 i24_4_lut_4_lut (.A(state[3]), .B(state[0]), .C(state[1]), .D(send), 
         .Z(n17)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i24_4_lut_4_lut.init = 16'h8001;
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n17_adj_299)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 i1_2_lut_rep_432 (.A(state[3]), .B(send), .Z(n28553)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_432.init = 16'h4444;
    LUT4 i20_4_lut_4_lut (.A(state[3]), .B(send), .C(state[0]), .D(state[1]), 
         .Z(n11)) /* synthesis lut_function=(A (C (D))+!A !((C+(D))+!B)) */ ;
    defparam i20_4_lut_4_lut.init = 16'ha004;
    LUT4 i2_3_lut (.A(\reset_count[7] ), .B(\reset_count[6] ), .C(\reset_count[5] ), 
         .Z(n24551)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i13_3_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), .D(state[3]), 
         .Z(n25937)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i13_3_lut_4_lut.init = 16'h0878;
    LUT4 i12_3_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), .D(state[3]), 
         .Z(n25763)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i12_3_lut_4_lut.init = 16'h0f80;
    LUT4 i20133_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n26829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20133_3_lut.init = 16'hcaca;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    LUT4 i8294_1_lut (.A(state[3]), .Z(n10070)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i8294_1_lut.init = 16'h5555;
    LUT4 i20134_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n26830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20134_3_lut.init = 16'hcaca;
    LUT4 i20316_4_lut_4_lut (.A(n28485), .B(n4), .C(n5020), .D(n1296), 
         .Z(n12642)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i20316_4_lut_4_lut.init = 16'h2a00;
    LUT4 i1_3_lut_3_lut (.A(n28485), .B(n11), .C(state[2]), .Z(n13549)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h5d5d;
    LUT4 i2_3_lut_3_lut (.A(n28485), .B(n1293), .C(n1290), .Z(n24779)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i2_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i2_4_lut (.A(n28553), .B(state[2]), .C(n19307), .D(n28485), 
         .Z(n8399)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0200;
    LUT4 i13329_2_lut (.A(state[1]), .B(state[0]), .Z(n19307)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13329_2_lut.init = 16'heeee;
    LUT4 i20447_3_lut (.A(n28485), .B(n17), .C(state[2]), .Z(n12687)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i20447_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut (.A(n28485), .B(state[1]), .C(n26766), .D(state[0]), 
         .Z(n26334)) /* synthesis lut_function=(!((B (C+(D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0208;
    LUT4 i20072_2_lut (.A(state[2]), .B(state[3]), .Z(n26766)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20072_2_lut.init = 16'h8888;
    FD1P3IX state__i2 (.D(n25937), .SP(n12687), .CD(n30473), .CK(bclk), 
            .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3IX state__i3 (.D(n25763), .SP(n12687), .CD(n30473), .CK(bclk), 
            .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1P3JX tx_35 (.D(n104), .SP(n17_adj_299), .PD(n30473), .CK(bclk), 
            .Q(n9969)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    FD1P3IX busy_34 (.D(n10070), .SP(n13549), .CD(n30473), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 state_2__bdd_4_lut_20731 (.A(state[0]), .B(state[3]), .C(state[1]), 
         .D(send), .Z(n27868)) /* synthesis lut_function=(A (B (C (D)))+!A (B+(C+(D)))) */ ;
    defparam state_2__bdd_4_lut_20731.init = 16'hd554;
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n26831), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i13479_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i13479_4_lut.init = 16'hfcee;
    \ClockDividerP(factor=12)  baud_gen (.GND_net(GND_net), .bclk(bclk), 
            .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (GND_net, bclk, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output bclk;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24360;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n102;
    
    wire n24359, n24358, n24357, n24356, n24355, n24354, n24353, 
        n24352, n55, n56, n4, n14871, n24351, n24060, n7556, 
        n24059, n24058, n52, n44, n24057, n24056, n24350, n35, 
        n54, n48, n36, n24349, n24348, n46, n32, n24055, n24054, 
        n24347, n50, n40, n24053, n24346, n24052, n24345, n24051, 
        n24050, n24049, n24048, n24047, n24046, n24045;
    
    CCU2D count_2377_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24360), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_33.INIT1 = 16'h0000;
    defparam count_2377_add_4_33.INJECT1_0 = "NO";
    defparam count_2377_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24359), .COUT(n24360), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_31.INJECT1_0 = "NO";
    defparam count_2377_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24358), .COUT(n24359), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_29.INJECT1_0 = "NO";
    defparam count_2377_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24357), .COUT(n24358), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_27.INJECT1_0 = "NO";
    defparam count_2377_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24356), .COUT(n24357), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_25.INJECT1_0 = "NO";
    defparam count_2377_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24355), .COUT(n24356), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_23.INJECT1_0 = "NO";
    defparam count_2377_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24354), .COUT(n24355), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_21.INJECT1_0 = "NO";
    defparam count_2377_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24353), .COUT(n24354), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_19.INJECT1_0 = "NO";
    defparam count_2377_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24352), .COUT(n24353), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_17.INJECT1_0 = "NO";
    defparam count_2377_add_4_17.INJECT1_1 = "NO";
    LUT4 i20353_4_lut (.A(n55), .B(count[1]), .C(n56), .D(n4), .Z(n14871)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20353_4_lut.init = 16'h0400;
    CCU2D count_2377_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24351), .COUT(n24352), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_15.INJECT1_0 = "NO";
    defparam count_2377_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24060), .S0(n7556));
    defparam sub_1888_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1888_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1888_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1888_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24059), .COUT(n24060));
    defparam sub_1888_add_2_32.INIT0 = 16'h5555;
    defparam sub_1888_add_2_32.INIT1 = 16'h5555;
    defparam sub_1888_add_2_32.INJECT1_0 = "NO";
    defparam sub_1888_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24058), .COUT(n24059));
    defparam sub_1888_add_2_30.INIT0 = 16'h5555;
    defparam sub_1888_add_2_30.INIT1 = 16'h5555;
    defparam sub_1888_add_2_30.INJECT1_0 = "NO";
    defparam sub_1888_add_2_30.INJECT1_1 = "NO";
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    CCU2D sub_1888_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24057), .COUT(n24058));
    defparam sub_1888_add_2_28.INIT0 = 16'h5555;
    defparam sub_1888_add_2_28.INIT1 = 16'h5555;
    defparam sub_1888_add_2_28.INJECT1_0 = "NO";
    defparam sub_1888_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24056), .COUT(n24057));
    defparam sub_1888_add_2_26.INIT0 = 16'h5555;
    defparam sub_1888_add_2_26.INIT1 = 16'h5555;
    defparam sub_1888_add_2_26.INJECT1_0 = "NO";
    defparam sub_1888_add_2_26.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24350), .COUT(n24351), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_13.INJECT1_0 = "NO";
    defparam count_2377_add_4_13.INJECT1_1 = "NO";
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[3]), .B(count[0]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    CCU2D count_2377_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24349), .COUT(n24350), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_11.INJECT1_0 = "NO";
    defparam count_2377_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24348), .COUT(n24349), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_9.INJECT1_0 = "NO";
    defparam count_2377_add_4_9.INJECT1_1 = "NO";
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    CCU2D sub_1888_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24055), .COUT(n24056));
    defparam sub_1888_add_2_24.INIT0 = 16'h5555;
    defparam sub_1888_add_2_24.INIT1 = 16'h5555;
    defparam sub_1888_add_2_24.INJECT1_0 = "NO";
    defparam sub_1888_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24054), .COUT(n24055));
    defparam sub_1888_add_2_22.INIT0 = 16'h5555;
    defparam sub_1888_add_2_22.INIT1 = 16'h5555;
    defparam sub_1888_add_2_22.INJECT1_0 = "NO";
    defparam sub_1888_add_2_22.INJECT1_1 = "NO";
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_3_lut.init = 16'hfefe;
    CCU2D count_2377_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24347), .COUT(n24348), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_7.INJECT1_0 = "NO";
    defparam count_2377_add_4_7.INJECT1_1 = "NO";
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i7_2_lut.init = 16'heeee;
    CCU2D sub_1888_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24053), .COUT(n24054));
    defparam sub_1888_add_2_20.INIT0 = 16'h5555;
    defparam sub_1888_add_2_20.INIT1 = 16'h5555;
    defparam sub_1888_add_2_20.INJECT1_0 = "NO";
    defparam sub_1888_add_2_20.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24346), .COUT(n24347), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_5.INJECT1_0 = "NO";
    defparam count_2377_add_4_5.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24052), .COUT(n24053));
    defparam sub_1888_add_2_18.INIT0 = 16'h5555;
    defparam sub_1888_add_2_18.INIT1 = 16'h5555;
    defparam sub_1888_add_2_18.INJECT1_0 = "NO";
    defparam sub_1888_add_2_18.INJECT1_1 = "NO";
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i11_2_lut.init = 16'heeee;
    CCU2D count_2377_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24345), .COUT(n24346), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2377_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2377_add_4_3.INJECT1_0 = "NO";
    defparam count_2377_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24051), .COUT(n24052));
    defparam sub_1888_add_2_16.INIT0 = 16'h5555;
    defparam sub_1888_add_2_16.INIT1 = 16'h5555;
    defparam sub_1888_add_2_16.INJECT1_0 = "NO";
    defparam sub_1888_add_2_16.INJECT1_1 = "NO";
    CCU2D count_2377_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24345), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377_add_4_1.INIT0 = 16'hF000;
    defparam count_2377_add_4_1.INIT1 = 16'h0555;
    defparam count_2377_add_4_1.INJECT1_0 = "NO";
    defparam count_2377_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24050), .COUT(n24051));
    defparam sub_1888_add_2_14.INIT0 = 16'h5555;
    defparam sub_1888_add_2_14.INIT1 = 16'h5555;
    defparam sub_1888_add_2_14.INJECT1_0 = "NO";
    defparam sub_1888_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24049), .COUT(n24050));
    defparam sub_1888_add_2_12.INIT0 = 16'h5555;
    defparam sub_1888_add_2_12.INIT1 = 16'h5555;
    defparam sub_1888_add_2_12.INJECT1_0 = "NO";
    defparam sub_1888_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24048), .COUT(n24049));
    defparam sub_1888_add_2_10.INIT0 = 16'h5555;
    defparam sub_1888_add_2_10.INIT1 = 16'h5555;
    defparam sub_1888_add_2_10.INJECT1_0 = "NO";
    defparam sub_1888_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24047), .COUT(n24048));
    defparam sub_1888_add_2_8.INIT0 = 16'h5555;
    defparam sub_1888_add_2_8.INIT1 = 16'h5555;
    defparam sub_1888_add_2_8.INJECT1_0 = "NO";
    defparam sub_1888_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24046), .COUT(n24047));
    defparam sub_1888_add_2_6.INIT0 = 16'h5555;
    defparam sub_1888_add_2_6.INIT1 = 16'h5555;
    defparam sub_1888_add_2_6.INJECT1_0 = "NO";
    defparam sub_1888_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24045), .COUT(n24046));
    defparam sub_1888_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1888_add_2_4.INIT1 = 16'h5555;
    defparam sub_1888_add_2_4.INJECT1_0 = "NO";
    defparam sub_1888_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_1888_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24045));
    defparam sub_1888_add_2_2.INIT0 = 16'h0000;
    defparam sub_1888_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1888_add_2_2.INJECT1_0 = "NO";
    defparam sub_1888_add_2_2.INJECT1_1 = "NO";
    FD1S3AX clk_o_14 (.D(n7556), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2377__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i0.GSR = "ENABLED";
    FD1S3IX count_2377__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i1.GSR = "ENABLED";
    FD1S3IX count_2377__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i2.GSR = "ENABLED";
    FD1S3IX count_2377__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i3.GSR = "ENABLED";
    FD1S3IX count_2377__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i4.GSR = "ENABLED";
    FD1S3IX count_2377__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i5.GSR = "ENABLED";
    FD1S3IX count_2377__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i6.GSR = "ENABLED";
    FD1S3IX count_2377__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i7.GSR = "ENABLED";
    FD1S3IX count_2377__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i8.GSR = "ENABLED";
    FD1S3IX count_2377__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i9.GSR = "ENABLED";
    FD1S3IX count_2377__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i10.GSR = "ENABLED";
    FD1S3IX count_2377__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i11.GSR = "ENABLED";
    FD1S3IX count_2377__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i12.GSR = "ENABLED";
    FD1S3IX count_2377__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i13.GSR = "ENABLED";
    FD1S3IX count_2377__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i14.GSR = "ENABLED";
    FD1S3IX count_2377__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i15.GSR = "ENABLED";
    FD1S3IX count_2377__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i16.GSR = "ENABLED";
    FD1S3IX count_2377__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i17.GSR = "ENABLED";
    FD1S3IX count_2377__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i18.GSR = "ENABLED";
    FD1S3IX count_2377__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i19.GSR = "ENABLED";
    FD1S3IX count_2377__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i20.GSR = "ENABLED";
    FD1S3IX count_2377__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i21.GSR = "ENABLED";
    FD1S3IX count_2377__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i22.GSR = "ENABLED";
    FD1S3IX count_2377__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i23.GSR = "ENABLED";
    FD1S3IX count_2377__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i24.GSR = "ENABLED";
    FD1S3IX count_2377__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i25.GSR = "ENABLED";
    FD1S3IX count_2377__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i26.GSR = "ENABLED";
    FD1S3IX count_2377__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i27.GSR = "ENABLED";
    FD1S3IX count_2377__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i28.GSR = "ENABLED";
    FD1S3IX count_2377__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i29.GSR = "ENABLED";
    FD1S3IX count_2377__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i30.GSR = "ENABLED";
    FD1S3IX count_2377__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n14871), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2377__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_c, n28485, rx_data, n30473, 
            n28457, debug_c_7, n9970_c, n28581, n28518, n28486, 
            n15, n12121, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n28485;
    output [7:0]rx_data;
    input n30473;
    input n28457;
    output debug_c_7;
    input n9970_c;
    output n28581;
    output n28518;
    output n28486;
    output n15;
    output n12121;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n8351, n8353;
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n25653, baud_reset, n19, n25221, n29248, n25351, n25579, 
        n25661, n8393, n8391, n8389, n8387, n8385, n8383, n8381, 
        n8379, n8377, n8375, n8373, n8371, n8369, n8367, n26580, 
        n25, n19_adj_294, n28469, n28590, n28589, bclk, n28549, 
        n19515, n10, n28501, n28556, n28559, n28470, n28557, n27, 
        n12356, n28558, n26586, n25_adj_295, n23, n26894, n21, 
        n23_adj_296, n12331, n19_adj_297;
    wire [7:0]n78;
    
    wire n13, n29247, n29245, n29246, n26616, n5, n27830, n28591, 
        n4, n9149, n4_adj_298, n26583;
    
    FD1P3AX rdata_i0_i0 (.D(n8351), .SP(n28485), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n8353), .SP(n28485), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n25653), .CK(debug_c_c), .CD(n30473), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n19), .CK(debug_c_c), .PD(n30473), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n25221), .CK(debug_c_c), .CD(n30473), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n29248), .CK(debug_c_c), .CD(n30473), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n25351), .CK(debug_c_c), .CD(n30473), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n25579), .CK(debug_c_c), .CD(n30473), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n25661), .CK(debug_c_c), .CD(n28457), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n8393), .SP(n28485), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n8391), .SP(n28485), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n8389), .SP(n28485), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n8387), .SP(n28485), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n8385), .SP(n28485), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n8383), .SP(n28485), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n8381), .SP(n28485), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n8379), .SP(n28485), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n8377), .SP(n28485), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n8375), .SP(n28485), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n8373), .SP(n28485), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n8371), .SP(n28485), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n8369), .SP(n28485), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i1 (.D(n8367), .SP(n28485), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    LUT4 i20373_4_lut (.A(debug_c_7), .B(n26580), .C(n9970_c), .D(n25), 
         .Z(n19_adj_294)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i20373_4_lut.init = 16'ha8ec;
    LUT4 i1_2_lut_rep_348_4_lut_4_lut (.A(state[4]), .B(state[3]), .C(state[2]), 
         .D(state[1]), .Z(n28469)) /* synthesis lut_function=(A+(B (C (D))+!B !(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_348_4_lut_4_lut.init = 16'heaab;
    LUT4 i1_3_lut_4_lut_4_lut_then_4_lut (.A(state[4]), .B(state[2]), .C(state[3]), 
         .D(state[1]), .Z(n28590)) /* synthesis lut_function=(A (C)+!A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_4_lut_then_4_lut.init = 16'he0a0;
    LUT4 i1_3_lut_4_lut_4_lut_else_4_lut (.A(state[4]), .B(state[2]), .C(state[3]), 
         .D(state[1]), .Z(n28589)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B !(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_4_lut_else_4_lut.init = 16'he0a1;
    LUT4 i13247_2_lut_rep_428 (.A(bclk), .B(state[1]), .Z(n28549)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13247_2_lut_rep_428.init = 16'h8888;
    LUT4 i13537_2_lut_3_lut (.A(bclk), .B(state[1]), .C(state[2]), .Z(n19515)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13537_2_lut_3_lut.init = 16'h8080;
    LUT4 i4_4_lut (.A(rx_data[3]), .B(rx_data[2]), .C(rx_data[1]), .D(rx_data[0]), 
         .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i4_4_lut.init = 16'h0100;
    LUT4 i1_3_lut_rep_380_4_lut (.A(state[2]), .B(state[1]), .C(state[3]), 
         .D(state[4]), .Z(n28501)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut_rep_380_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_435 (.A(state[1]), .B(state[4]), .Z(n28556)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_435.init = 16'heeee;
    LUT4 i19980_2_lut_rep_349_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(n9970_c), 
         .D(n28559), .Z(n28470)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i19980_2_lut_rep_349_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(n28557), 
         .D(n28559), .Z(n26580)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_173 (.A(state[1]), .B(state[4]), .C(n28559), 
         .D(state[0]), .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut_adj_173.init = 16'hfffe;
    LUT4 i41_4_lut_3_lut (.A(bclk), .B(state[1]), .C(state[2]), .Z(n27)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i41_4_lut_3_lut.init = 16'hb4b4;
    LUT4 i13008_2_lut_rep_436 (.A(state[0]), .B(state[5]), .Z(n28557)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13008_2_lut_rep_436.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n12356)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_437 (.A(state[1]), .B(bclk), .Z(n28558)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_rep_437.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_174 (.A(state[1]), .B(bclk), .C(state[2]), 
         .Z(n26586)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_3_lut_adj_174.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_438 (.A(state[2]), .B(state[3]), .Z(n28559)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_rep_438.init = 16'heeee;
    FD1S3IX drdy_51 (.D(n19_adj_294), .CK(debug_c_c), .CD(n30473), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    PFUMX i40 (.BLUT(n25_adj_295), .ALUT(n27), .C0(state[0]), .Z(n25579));
    PFUMX i36 (.BLUT(n23), .ALUT(n26894), .C0(state[0]), .Z(n25661));
    PFUMX i36_adj_175 (.BLUT(n21), .ALUT(n23_adj_296), .C0(state[5]), 
          .Z(n25221));
    LUT4 i2_3_lut_4_lut (.A(n28559), .B(n28556), .C(state[0]), .D(state[5]), 
         .Z(n12331)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_4_lut_adj_176 (.A(state[0]), .B(n28556), .C(state[5]), 
         .D(n28559), .Z(n19_adj_297)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_4_lut_adj_176.init = 16'hffef;
    LUT4 i1_4_lut (.A(n78[0]), .B(rdata[0]), .C(n12356), .D(n13), .Z(n8351)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i4100_4_lut (.A(n9970_c), .B(rdata[0]), .C(n28559), .D(n28558), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4100_4_lut.init = 16'hccca;
    LUT4 i32_2_lut_rep_460 (.A(rx_data[6]), .B(rx_data[7]), .Z(n28581)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i32_2_lut_rep_460.init = 16'heeee;
    LUT4 i20096_2_lut_rep_397_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(rx_data[5]), 
         .Z(n28518)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i20096_2_lut_rep_397_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut.init = 16'hefef;
    LUT4 state_4__bdd_2_lut (.A(state[4]), .B(state[5]), .Z(n29247)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam state_4__bdd_2_lut.init = 16'h2222;
    LUT4 state_4__bdd_3_lut (.A(state[4]), .B(n29245), .C(state[2]), .Z(n29246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam state_4__bdd_3_lut.init = 16'hcaca;
    LUT4 state_4__bdd_4_lut_21314 (.A(state[4]), .B(bclk), .C(state[3]), 
         .D(state[1]), .Z(n29245)) /* synthesis lut_function=(A (B+!(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam state_4__bdd_4_lut_21314.init = 16'h9aaa;
    LUT4 i5_3_lut_rep_365_4_lut (.A(rx_data[5]), .B(n28581), .C(rx_data[4]), 
         .D(n10), .Z(n28486)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i5_3_lut_rep_365_4_lut.init = 16'h0100;
    LUT4 i3_4_lut (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), .D(n26616), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n26616), .B(rx_data[4]), .C(rx_data[1]), .D(rx_data[3]), 
         .Z(n12121)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'hbfff;
    LUT4 i1_4_lut_adj_177 (.A(rx_data[2]), .B(n5), .C(rx_data[0]), .D(rx_data[7]), 
         .Z(n26616)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_177.init = 16'hffef;
    LUT4 i1_2_lut (.A(rx_data[5]), .B(rx_data[6]), .Z(n5)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_178 (.A(rdata[0]), .B(rx_data[0]), .C(n12331), .D(n19_adj_297), 
         .Z(n8353)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_178.init = 16'heca0;
    LUT4 i1_4_lut_adj_179 (.A(state[5]), .B(n28470), .C(state[2]), .D(n28469), 
         .Z(n25_adj_295)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_179.init = 16'h5111;
    LUT4 i20375_4_lut (.A(baud_reset), .B(n26580), .C(n9970_c), .D(n25), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i20375_4_lut.init = 16'ha8ec;
    LUT4 i1_4_lut_adj_180 (.A(state[5]), .B(n28470), .C(state[1]), .D(n28469), 
         .Z(n23)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_180.init = 16'h5111;
    LUT4 i20295_2_lut (.A(bclk), .B(state[1]), .Z(n26894)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i20295_2_lut.init = 16'h9999;
    LUT4 i43_4_lut (.A(state[5]), .B(n27830), .C(state[0]), .D(n28591), 
         .Z(n25351)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i43_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_adj_181 (.A(rdata[7]), .B(rx_data[7]), .C(n12331), .D(n19_adj_297), 
         .Z(n8393)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_181.init = 16'heca0;
    LUT4 i1_4_lut_adj_182 (.A(rdata[6]), .B(rx_data[6]), .C(n12331), .D(n19_adj_297), 
         .Z(n8391)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_182.init = 16'heca0;
    LUT4 i1_4_lut_adj_183 (.A(rdata[5]), .B(rx_data[5]), .C(n12331), .D(n19_adj_297), 
         .Z(n8389)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_183.init = 16'heca0;
    LUT4 i1_4_lut_adj_184 (.A(rdata[4]), .B(rx_data[4]), .C(n12331), .D(n19_adj_297), 
         .Z(n8387)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_184.init = 16'heca0;
    LUT4 i2_4_lut_adj_185 (.A(bclk), .B(n4), .C(state[0]), .D(n28501), 
         .Z(n21)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut_adj_185.init = 16'h4840;
    LUT4 i1_2_lut_adj_186 (.A(state[4]), .B(n9149), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_186.init = 16'h8888;
    LUT4 i38_4_lut (.A(n28470), .B(n9149), .C(state[0]), .D(n4_adj_298), 
         .Z(n23_adj_296)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i38_4_lut.init = 16'hf535;
    LUT4 i1_2_lut_adj_187 (.A(state[4]), .B(bclk), .Z(n4_adj_298)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_187.init = 16'hdddd;
    LUT4 i1_4_lut_adj_188 (.A(rdata[3]), .B(rx_data[3]), .C(n12331), .D(n19_adj_297), 
         .Z(n8385)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_188.init = 16'heca0;
    LUT4 i1_4_lut_adj_189 (.A(rdata[2]), .B(rx_data[2]), .C(n12331), .D(n19_adj_297), 
         .Z(n8383)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_189.init = 16'heca0;
    LUT4 i1_4_lut_adj_190 (.A(rdata[1]), .B(rx_data[1]), .C(n12331), .D(n19_adj_297), 
         .Z(n8381)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_190.init = 16'heca0;
    LUT4 i3123_4_lut (.A(state[3]), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(n9149)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3123_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_191 (.A(n78[7]), .B(rdata[7]), .C(n12356), .D(n13), 
         .Z(n8379)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_191.init = 16'heca0;
    LUT4 i4040_4_lut (.A(rdata[7]), .B(n9970_c), .C(state[3]), .D(n19515), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4040_4_lut.init = 16'hcaaa;
    LUT4 i1_4_lut_adj_192 (.A(n78[6]), .B(rdata[6]), .C(n12356), .D(n13), 
         .Z(n8377)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_192.init = 16'heca0;
    LUT4 i4042_4_lut (.A(n9970_c), .B(rdata[6]), .C(state[3]), .D(n26586), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4042_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_193 (.A(n78[5]), .B(rdata[5]), .C(n12356), .D(n13), 
         .Z(n8375)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_193.init = 16'heca0;
    LUT4 i4044_4_lut (.A(n9970_c), .B(rdata[5]), .C(n28549), .D(n26583), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4044_4_lut.init = 16'hccac;
    LUT4 i1_2_lut_adj_194 (.A(state[2]), .B(state[3]), .Z(n26583)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_adj_194.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_195 (.A(n78[4]), .B(rdata[4]), .C(n12356), .D(n13), 
         .Z(n8373)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_195.init = 16'heca0;
    LUT4 i4046_4_lut (.A(n9970_c), .B(rdata[4]), .C(n28558), .D(n26583), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4046_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_196 (.A(n78[3]), .B(rdata[3]), .C(n12356), .D(n13), 
         .Z(n8371)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_196.init = 16'heca0;
    LUT4 i4048_4_lut (.A(n9970_c), .B(rdata[3]), .C(state[3]), .D(n19515), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4048_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_197 (.A(n78[2]), .B(rdata[2]), .C(n12356), .D(n13), 
         .Z(n8369)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_197.init = 16'heca0;
    LUT4 i4050_4_lut (.A(n9970_c), .B(rdata[2]), .C(state[3]), .D(n26586), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4050_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_198 (.A(n78[1]), .B(rdata[1]), .C(n12356), .D(n13), 
         .Z(n8367)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_198.init = 16'heca0;
    LUT4 i4052_4_lut (.A(n9970_c), .B(rdata[1]), .C(n28559), .D(n28549), 
         .Z(n78[1])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4052_4_lut.init = 16'hcacc;
    PFUMX i21220 (.BLUT(n29247), .ALUT(n29246), .C0(state[0]), .Z(n29248));
    LUT4 state_3__bdd_4_lut_21241 (.A(state[3]), .B(bclk), .C(state[2]), 
         .D(state[1]), .Z(n27830)) /* synthesis lut_function=(A (B+!(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam state_3__bdd_4_lut_21241.init = 16'h9aaa;
    LUT4 i1_3_lut_4_lut (.A(state[5]), .B(n28501), .C(state[0]), .D(bclk), 
         .Z(n25653)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut.init = 16'hf400;
    PFUMX i20880 (.BLUT(n28589), .ALUT(n28590), .C0(n9970_c), .Z(n28591));
    \ClockDividerP(factor=12)_U0  baud_gen (.GND_net(GND_net), .bclk(bclk), 
            .debug_c_c(debug_c_c), .baud_reset(baud_reset)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (GND_net, bclk, debug_c_c, baud_reset) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output bclk;
    input debug_c_c;
    input baud_reset;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n24409, n7521, n2732;
    wire [31:0]n134;
    
    wire n24312, n24311, n24310, n24309, n24308, n24307, n24306, 
        n24305, n24304, n24303, n24302, n24301, n24300, n24299, 
        n24298, n24297, n55, n24622, n56, n52, n44, n35, n54, 
        n48, n36, n46, n32, n50, n40, n24424, n24423, n24422, 
        n24421, n24420, n24419, n24418, n24417, n24416, n24415, 
        n24414, n24413, n24412, n24411, n24410;
    
    CCU2D sub_1886_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24409));
    defparam sub_1886_add_2_2.INIT0 = 16'h0000;
    defparam sub_1886_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1886_add_2_2.INJECT1_0 = "NO";
    defparam sub_1886_add_2_2.INJECT1_1 = "NO";
    FD1S3IX clk_o_14 (.D(n7521), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2376__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2732), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i0.GSR = "ENABLED";
    CCU2D count_2376_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24312), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_33.INIT1 = 16'h0000;
    defparam count_2376_add_4_33.INJECT1_0 = "NO";
    defparam count_2376_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24311), .COUT(n24312), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_31.INJECT1_0 = "NO";
    defparam count_2376_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24310), .COUT(n24311), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_29.INJECT1_0 = "NO";
    defparam count_2376_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24309), .COUT(n24310), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_27.INJECT1_0 = "NO";
    defparam count_2376_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24308), .COUT(n24309), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_25.INJECT1_0 = "NO";
    defparam count_2376_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24307), .COUT(n24308), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_23.INJECT1_0 = "NO";
    defparam count_2376_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24306), .COUT(n24307), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_21.INJECT1_0 = "NO";
    defparam count_2376_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24305), .COUT(n24306), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_19.INJECT1_0 = "NO";
    defparam count_2376_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24304), .COUT(n24305), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_17.INJECT1_0 = "NO";
    defparam count_2376_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24303), .COUT(n24304), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_15.INJECT1_0 = "NO";
    defparam count_2376_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24302), .COUT(n24303), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_13.INJECT1_0 = "NO";
    defparam count_2376_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24301), .COUT(n24302), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_11.INJECT1_0 = "NO";
    defparam count_2376_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24300), .COUT(n24301), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_9.INJECT1_0 = "NO";
    defparam count_2376_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24299), .COUT(n24300), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_7.INJECT1_0 = "NO";
    defparam count_2376_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24298), .COUT(n24299), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_5.INJECT1_0 = "NO";
    defparam count_2376_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24297), .COUT(n24298), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2376_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2376_add_4_3.INJECT1_0 = "NO";
    defparam count_2376_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2376_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24297), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376_add_4_1.INIT0 = 16'hF000;
    defparam count_2376_add_4_1.INIT1 = 16'h0555;
    defparam count_2376_add_4_1.INJECT1_0 = "NO";
    defparam count_2376_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2376__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2732), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i1.GSR = "ENABLED";
    FD1S3IX count_2376__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2732), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i2.GSR = "ENABLED";
    FD1S3IX count_2376__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2732), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i3.GSR = "ENABLED";
    FD1S3IX count_2376__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2732), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i4.GSR = "ENABLED";
    FD1S3IX count_2376__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2732), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i5.GSR = "ENABLED";
    FD1S3IX count_2376__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2732), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i6.GSR = "ENABLED";
    FD1S3IX count_2376__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2732), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i7.GSR = "ENABLED";
    FD1S3IX count_2376__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2732), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i8.GSR = "ENABLED";
    FD1S3IX count_2376__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2732), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i9.GSR = "ENABLED";
    FD1S3IX count_2376__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i10.GSR = "ENABLED";
    FD1S3IX count_2376__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i11.GSR = "ENABLED";
    FD1S3IX count_2376__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i12.GSR = "ENABLED";
    FD1S3IX count_2376__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i13.GSR = "ENABLED";
    FD1S3IX count_2376__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i14.GSR = "ENABLED";
    FD1S3IX count_2376__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i15.GSR = "ENABLED";
    FD1S3IX count_2376__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i16.GSR = "ENABLED";
    FD1S3IX count_2376__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i17.GSR = "ENABLED";
    FD1S3IX count_2376__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i18.GSR = "ENABLED";
    FD1S3IX count_2376__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i19.GSR = "ENABLED";
    FD1S3IX count_2376__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i20.GSR = "ENABLED";
    FD1S3IX count_2376__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i21.GSR = "ENABLED";
    FD1S3IX count_2376__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i22.GSR = "ENABLED";
    FD1S3IX count_2376__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i23.GSR = "ENABLED";
    FD1S3IX count_2376__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i24.GSR = "ENABLED";
    FD1S3IX count_2376__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i25.GSR = "ENABLED";
    FD1S3IX count_2376__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i26.GSR = "ENABLED";
    FD1S3IX count_2376__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i27.GSR = "ENABLED";
    FD1S3IX count_2376__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i28.GSR = "ENABLED";
    FD1S3IX count_2376__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i29.GSR = "ENABLED";
    FD1S3IX count_2376__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i30.GSR = "ENABLED";
    FD1S3IX count_2376__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2732), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2376__i31.GSR = "ENABLED";
    LUT4 i1056_4_lut (.A(n55), .B(baud_reset), .C(n24622), .D(n56), 
         .Z(n2732)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i1056_4_lut.init = 16'hccdc;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(count[1]), .B(count[3]), .C(count[0]), .Z(n24622)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_2_lut.init = 16'heeee;
    CCU2D sub_1886_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24424), .S0(n7521));
    defparam sub_1886_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1886_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1886_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1886_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24423), .COUT(n24424));
    defparam sub_1886_add_2_32.INIT0 = 16'h5555;
    defparam sub_1886_add_2_32.INIT1 = 16'h5555;
    defparam sub_1886_add_2_32.INJECT1_0 = "NO";
    defparam sub_1886_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24422), .COUT(n24423));
    defparam sub_1886_add_2_30.INIT0 = 16'h5555;
    defparam sub_1886_add_2_30.INIT1 = 16'h5555;
    defparam sub_1886_add_2_30.INJECT1_0 = "NO";
    defparam sub_1886_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24421), .COUT(n24422));
    defparam sub_1886_add_2_28.INIT0 = 16'h5555;
    defparam sub_1886_add_2_28.INIT1 = 16'h5555;
    defparam sub_1886_add_2_28.INJECT1_0 = "NO";
    defparam sub_1886_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24420), .COUT(n24421));
    defparam sub_1886_add_2_26.INIT0 = 16'h5555;
    defparam sub_1886_add_2_26.INIT1 = 16'h5555;
    defparam sub_1886_add_2_26.INJECT1_0 = "NO";
    defparam sub_1886_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24419), .COUT(n24420));
    defparam sub_1886_add_2_24.INIT0 = 16'h5555;
    defparam sub_1886_add_2_24.INIT1 = 16'h5555;
    defparam sub_1886_add_2_24.INJECT1_0 = "NO";
    defparam sub_1886_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24418), .COUT(n24419));
    defparam sub_1886_add_2_22.INIT0 = 16'h5555;
    defparam sub_1886_add_2_22.INIT1 = 16'h5555;
    defparam sub_1886_add_2_22.INJECT1_0 = "NO";
    defparam sub_1886_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24417), .COUT(n24418));
    defparam sub_1886_add_2_20.INIT0 = 16'h5555;
    defparam sub_1886_add_2_20.INIT1 = 16'h5555;
    defparam sub_1886_add_2_20.INJECT1_0 = "NO";
    defparam sub_1886_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24416), .COUT(n24417));
    defparam sub_1886_add_2_18.INIT0 = 16'h5555;
    defparam sub_1886_add_2_18.INIT1 = 16'h5555;
    defparam sub_1886_add_2_18.INJECT1_0 = "NO";
    defparam sub_1886_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24415), .COUT(n24416));
    defparam sub_1886_add_2_16.INIT0 = 16'h5555;
    defparam sub_1886_add_2_16.INIT1 = 16'h5555;
    defparam sub_1886_add_2_16.INJECT1_0 = "NO";
    defparam sub_1886_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24414), .COUT(n24415));
    defparam sub_1886_add_2_14.INIT0 = 16'h5555;
    defparam sub_1886_add_2_14.INIT1 = 16'h5555;
    defparam sub_1886_add_2_14.INJECT1_0 = "NO";
    defparam sub_1886_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24413), .COUT(n24414));
    defparam sub_1886_add_2_12.INIT0 = 16'h5555;
    defparam sub_1886_add_2_12.INIT1 = 16'h5555;
    defparam sub_1886_add_2_12.INJECT1_0 = "NO";
    defparam sub_1886_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24412), .COUT(n24413));
    defparam sub_1886_add_2_10.INIT0 = 16'h5555;
    defparam sub_1886_add_2_10.INIT1 = 16'h5555;
    defparam sub_1886_add_2_10.INJECT1_0 = "NO";
    defparam sub_1886_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24411), .COUT(n24412));
    defparam sub_1886_add_2_8.INIT0 = 16'h5555;
    defparam sub_1886_add_2_8.INIT1 = 16'h5555;
    defparam sub_1886_add_2_8.INJECT1_0 = "NO";
    defparam sub_1886_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24410), .COUT(n24411));
    defparam sub_1886_add_2_6.INIT0 = 16'h5555;
    defparam sub_1886_add_2_6.INIT1 = 16'h5555;
    defparam sub_1886_add_2_6.INJECT1_0 = "NO";
    defparam sub_1886_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1886_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24409), .COUT(n24410));
    defparam sub_1886_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1886_add_2_4.INIT1 = 16'h5555;
    defparam sub_1886_add_2_4.INJECT1_0 = "NO";
    defparam sub_1886_add_2_4.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (\register_addr[0] , \register_addr[2] , \register_addr[1] , 
            \select[7] , n176, databus_out, n2, rw, databus, \read_value[12] , 
            n1, n28582, \read_value[12]_adj_6 , read_value, n28451, 
            n52, n2_adj_8, n2_adj_9, n2_adj_10, \read_value[8]_adj_11 , 
            n1_adj_12, \read_value[8]_adj_13 , \read_value[9]_adj_14 , 
            n1_adj_15, read_size, \read_size[0]_adj_16 , \select[1] , 
            n28487, n9, \read_size[0]_adj_17 , n28452, n28476, \read_size[0]_adj_18 , 
            n10, \read_size[0]_adj_19 , \select[2] , n8, \read_size[2]_adj_20 , 
            \reg_size[2] , \read_size[2]_adj_21 , \read_size[2]_adj_22 , 
            \read_size[2]_adj_23 , n28480, n4, \read_value[0]_adj_24 , 
            n28448, \read_value[0]_adj_25 , \read_value[0]_adj_26 , n28458, 
            read_value_adj_146, n64, n2_adj_35, \read_value[9]_adj_36 , 
            n2_adj_37, \read_value[21]_adj_38 , n1_adj_39, \read_value[31]_adj_40 , 
            n1_adj_41, \read_value[31]_adj_42 , n4_adj_43, \read_value[7]_adj_44 , 
            n28576, \sendcount[1] , n11943, n28439, \read_value[13]_adj_45 , 
            n1_adj_46, n4_adj_47, \read_value[6]_adj_48 , \read_value[7]_adj_49 , 
            \read_value[7]_adj_50 , \read_value[13]_adj_51 , \read_value[6]_adj_52 , 
            \read_value[6]_adj_53 , n2_adj_54, \read_value[21]_adj_55 , 
            \read_value[11]_adj_56 , n1_adj_57, \read_value[10]_adj_58 , 
            n2_adj_59, \read_value[30]_adj_60 , n1_adj_61, n4_adj_62, 
            \read_value[5]_adj_63 , \read_value[5]_adj_64 , \read_value[5]_adj_65 , 
            n30468, \read_value[30]_adj_66 , n4_adj_67, \read_value[4]_adj_68 , 
            \read_value[4]_adj_69 , \read_value[4]_adj_70 , n4_adj_71, 
            \read_value[2]_adj_72 , \read_value[2]_adj_73 , \read_value[2]_adj_74 , 
            \read_value[11]_adj_75 , n2_adj_76, \read_value[28]_adj_77 , 
            n1_adj_78, \read_value[28]_adj_79 , n2_adj_80, \read_value[27]_adj_81 , 
            n1_adj_82, n1_adj_83, n2_adj_84, \read_value[1]_adj_85 , 
            n6, n2_adj_86, \read_value[20]_adj_87 , n1_adj_88, \read_value[27]_adj_89 , 
            n2_adj_90, \read_value[20]_adj_91 , n2_adj_92, \read_value[14]_adj_93 , 
            n1_adj_94, \read_value[14]_adj_95 , \read_value[19]_adj_96 , 
            n1_adj_97, n4_adj_98, \read_value[10]_adj_99 , n1_adj_100, 
            \read_value[3]_adj_101 , n2_adj_102, \read_value[19]_adj_103 , 
            \read_value[26]_adj_104 , n1_adj_105, \read_value[3]_adj_106 , 
            \read_value[3]_adj_107 , \read_value[26]_adj_108 , n2_adj_109, 
            \read_value[25]_adj_110 , n1_adj_111, n2_adj_112, \read_value[18]_adj_113 , 
            n1_adj_114, \read_value[25]_adj_115 , \read_value[18]_adj_116 , 
            n2_adj_117, \read_value[17]_adj_118 , n1_adj_119, \read_value[17]_adj_120 , 
            n2_adj_121, \read_value[24]_adj_122 , n1_adj_123, \read_value[24]_adj_124 , 
            \read_value[1]_adj_125 , n2_adj_126, \read_value[16]_adj_127 , 
            n1_adj_128, n2_adj_129, n2_adj_130, \read_value[29]_adj_131 , 
            n1_adj_132, \read_value[16]_adj_133 , \read_value[29]_adj_134 , 
            \read_value[23]_adj_135 , n1_adj_136, n2_adj_137, \read_value[23]_adj_138 , 
            \read_value[15]_adj_139 , n1_adj_140, n2_adj_141, \read_value[22]_adj_142 , 
            n1_adj_143, \read_value[15]_adj_144 , \read_value[22]_adj_145 , 
            debug_c_c, n30470, rc_ch8_c, GND_net, n26922, n30469, 
            n26942, n12605, n24743, n30471, n13489, rc_ch7_c, n26949, 
            n24707, n27040, n13527, rc_ch4_c, n26947, n24721, n27035, 
            n13534, rc_ch3_c, n27027, n26939, n24755, rc_ch2_c, 
            n26945, n13535, n24741, n27025, n28403, n26907, rc_ch1_c, 
            n13536, n24716, n27023) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[0] ;
    input \register_addr[2] ;
    input \register_addr[1] ;
    input \select[7] ;
    input n176;
    input [31:0]databus_out;
    input n2;
    input rw;
    output [31:0]databus;
    input \read_value[12] ;
    input n1;
    input n28582;
    input \read_value[12]_adj_6 ;
    input [31:0]read_value;
    input n28451;
    input n52;
    input n2_adj_8;
    input n2_adj_9;
    input n2_adj_10;
    input \read_value[8]_adj_11 ;
    input n1_adj_12;
    input \read_value[8]_adj_13 ;
    input \read_value[9]_adj_14 ;
    input n1_adj_15;
    input [2:0]read_size;
    input \read_size[0]_adj_16 ;
    input \select[1] ;
    input n28487;
    output n9;
    input \read_size[0]_adj_17 ;
    input n28452;
    input n28476;
    input \read_size[0]_adj_18 ;
    output n10;
    input \read_size[0]_adj_19 ;
    input \select[2] ;
    output n8;
    input \read_size[2]_adj_20 ;
    output \reg_size[2] ;
    input \read_size[2]_adj_21 ;
    input \read_size[2]_adj_22 ;
    input \read_size[2]_adj_23 ;
    input n28480;
    input n4;
    input \read_value[0]_adj_24 ;
    input n28448;
    input \read_value[0]_adj_25 ;
    input \read_value[0]_adj_26 ;
    input n28458;
    input [7:0]read_value_adj_146;
    input n64;
    input n2_adj_35;
    input \read_value[9]_adj_36 ;
    input n2_adj_37;
    input \read_value[21]_adj_38 ;
    input n1_adj_39;
    input \read_value[31]_adj_40 ;
    input n1_adj_41;
    input \read_value[31]_adj_42 ;
    input n4_adj_43;
    input \read_value[7]_adj_44 ;
    output n28576;
    input \sendcount[1] ;
    output n11943;
    input n28439;
    input \read_value[13]_adj_45 ;
    input n1_adj_46;
    input n4_adj_47;
    input \read_value[6]_adj_48 ;
    input \read_value[7]_adj_49 ;
    input \read_value[7]_adj_50 ;
    input \read_value[13]_adj_51 ;
    input \read_value[6]_adj_52 ;
    input \read_value[6]_adj_53 ;
    input n2_adj_54;
    input \read_value[21]_adj_55 ;
    input \read_value[11]_adj_56 ;
    input n1_adj_57;
    input \read_value[10]_adj_58 ;
    input n2_adj_59;
    input \read_value[30]_adj_60 ;
    input n1_adj_61;
    input n4_adj_62;
    input \read_value[5]_adj_63 ;
    input \read_value[5]_adj_64 ;
    input \read_value[5]_adj_65 ;
    input n30468;
    input \read_value[30]_adj_66 ;
    input n4_adj_67;
    input \read_value[4]_adj_68 ;
    input \read_value[4]_adj_69 ;
    input \read_value[4]_adj_70 ;
    input n4_adj_71;
    input \read_value[2]_adj_72 ;
    input \read_value[2]_adj_73 ;
    input \read_value[2]_adj_74 ;
    input \read_value[11]_adj_75 ;
    input n2_adj_76;
    input \read_value[28]_adj_77 ;
    input n1_adj_78;
    input \read_value[28]_adj_79 ;
    input n2_adj_80;
    input \read_value[27]_adj_81 ;
    input n1_adj_82;
    input n1_adj_83;
    input n2_adj_84;
    input \read_value[1]_adj_85 ;
    input n6;
    input n2_adj_86;
    input \read_value[20]_adj_87 ;
    input n1_adj_88;
    input \read_value[27]_adj_89 ;
    input n2_adj_90;
    input \read_value[20]_adj_91 ;
    input n2_adj_92;
    input \read_value[14]_adj_93 ;
    input n1_adj_94;
    input \read_value[14]_adj_95 ;
    input \read_value[19]_adj_96 ;
    input n1_adj_97;
    input n4_adj_98;
    input \read_value[10]_adj_99 ;
    input n1_adj_100;
    input \read_value[3]_adj_101 ;
    input n2_adj_102;
    input \read_value[19]_adj_103 ;
    input \read_value[26]_adj_104 ;
    input n1_adj_105;
    input \read_value[3]_adj_106 ;
    input \read_value[3]_adj_107 ;
    input \read_value[26]_adj_108 ;
    input n2_adj_109;
    input \read_value[25]_adj_110 ;
    input n1_adj_111;
    input n2_adj_112;
    input \read_value[18]_adj_113 ;
    input n1_adj_114;
    input \read_value[25]_adj_115 ;
    input \read_value[18]_adj_116 ;
    input n2_adj_117;
    input \read_value[17]_adj_118 ;
    input n1_adj_119;
    input \read_value[17]_adj_120 ;
    input n2_adj_121;
    input \read_value[24]_adj_122 ;
    input n1_adj_123;
    input \read_value[24]_adj_124 ;
    input \read_value[1]_adj_125 ;
    input n2_adj_126;
    input \read_value[16]_adj_127 ;
    input n1_adj_128;
    input n2_adj_129;
    input n2_adj_130;
    input \read_value[29]_adj_131 ;
    input n1_adj_132;
    input \read_value[16]_adj_133 ;
    input \read_value[29]_adj_134 ;
    input \read_value[23]_adj_135 ;
    input n1_adj_136;
    input n2_adj_137;
    input \read_value[23]_adj_138 ;
    input \read_value[15]_adj_139 ;
    input n1_adj_140;
    input n2_adj_141;
    input \read_value[22]_adj_142 ;
    input n1_adj_143;
    input \read_value[15]_adj_144 ;
    input \read_value[22]_adj_145 ;
    input debug_c_c;
    input n30470;
    input rc_ch8_c;
    input GND_net;
    output n26922;
    input n30469;
    output n26942;
    input n12605;
    input n24743;
    input n30471;
    input n13489;
    input rc_ch7_c;
    output n26949;
    input n24707;
    output n27040;
    input n13527;
    input rc_ch4_c;
    output n26947;
    input n24721;
    output n27035;
    input n13534;
    input rc_ch3_c;
    output n27027;
    output n26939;
    input n24755;
    input rc_ch2_c;
    output n26945;
    input n13535;
    input n24741;
    output n27025;
    input n28403;
    output n26907;
    input rc_ch1_c;
    input n13536;
    input n24716;
    output n27023;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n971;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n27692;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n27691;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n27688, n28381;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n28382, n27828, n27825, n27829, n27827, n27826, n28384;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(211[12:21])
    
    wire n1031, n28385, n27824, n27823, n27812, n27809, n27813, 
        n27811, n27810, n27808, n27807, n27405, n27406, n10_c, 
        n8_c, n27408, n1016, n27409, n986, n27464, n27994, n27992, 
        n27991, n27995, n10_adj_59, n10_adj_61, n10_adj_63, n8_adj_65, 
        n8_adj_69, n7, n6_c, n28568;
    wire [7:0]read_value_adj_292;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(210[12:22])
    
    wire n7_adj_82, n7_adj_83, n7_adj_84, n7_adj_85, n7_adj_86, n7_adj_87, 
        n7_adj_88, n13, n12, n6_adj_89, n10_adj_91, n10_adj_96, 
        n28233, n10_adj_100, n8_adj_102, n8_adj_104, n28232, n28235, 
        n28236, n13_adj_108, n12_adj_110, n6_adj_111, n27465, n27462, 
        n27466, n10_adj_113, n28387, n28238, n27997, n27411, n8_adj_114, 
        n13_adj_116, n12_adj_118, n6_adj_119, n10_adj_121, n10_adj_128, 
        n27463, n27689, n8_adj_136, n8_adj_139, n27461, n27460, 
        n1001, n10_adj_140, n8_adj_142, n13_adj_144, n12_adj_146, 
        n6_adj_147, n10_adj_149, n27410, n27407, n13_adj_156, n12_adj_158, 
        n6_adj_159, n10_adj_161, n27693, n27690, n27694, n13_adj_166, 
        n12_adj_168, n6_adj_169, n10_adj_171, n28386, n28383, n1046, 
        n10_adj_178, n8_adj_180, n10_adj_184, n8_adj_186, n14, n10_adj_189, 
        n7_adj_190, n10_adj_191, n12_adj_194, n10_adj_196, n8_adj_198, 
        n10_adj_202, n10_adj_206, n8_adj_208, n28237, n28234, n8_adj_214, 
        n13_adj_216, n12_adj_218, n6_adj_219, n10_adj_223, n10_adj_224, 
        n8_adj_228, n10_adj_234, n8_adj_236, n10_adj_238, n8_adj_240, 
        n10_adj_248, n8_adj_250, n10_adj_254, n27996, n27993, n8_adj_256, 
        n10_adj_261, n8_adj_263, n10_adj_265, n10_adj_267, n8_adj_269, 
        n8_adj_275, n10_adj_277, n8_adj_281, n10_adj_283, n8_adj_285;
    
    LUT4 n971_bdd_3_lut_20695 (.A(n971), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n27692)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n971_bdd_3_lut_20695.init = 16'he2e2;
    LUT4 n971_bdd_3_lut_20614 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n27691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n971_bdd_3_lut_20614.init = 16'hcaca;
    LUT4 register_addr_1__bdd_2_lut_20659 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n27688)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_20659.init = 16'h2222;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n28381)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n28382)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    L6MUX21 i20680 (.D0(n27828), .D1(n27825), .SD(\register_addr[2] ), 
            .Z(n27829));
    PFUMX i20678 (.BLUT(n27827), .ALUT(n27826), .C0(\register_addr[1] ), 
          .Z(n27828));
    LUT4 n1031_bdd_3_lut_20865 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n28384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1031_bdd_3_lut_20865.init = 16'hcaca;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 n1031_bdd_3_lut_21294 (.A(n1031), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n28385)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1031_bdd_3_lut_21294.init = 16'he2e2;
    PFUMX i20675 (.BLUT(n27824), .ALUT(n27823), .C0(\register_addr[1] ), 
          .Z(n27825));
    L6MUX21 i20668 (.D0(n27812), .D1(n27809), .SD(\register_addr[2] ), 
            .Z(n27813));
    LUT4 n1046_bdd_3_lut_20677 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n27826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1046_bdd_3_lut_20677.init = 16'hcaca;
    PFUMX i20666 (.BLUT(n27811), .ALUT(n27810), .C0(\register_addr[1] ), 
          .Z(n27812));
    PFUMX i20663 (.BLUT(n27808), .ALUT(n27807), .C0(\register_addr[1] ), 
          .Z(n27809));
    LUT4 register_addr_1__bdd_2_lut_20545 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n27405)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_20545.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_20546 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n27406)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_20546.init = 16'he4e4;
    LUT4 i5_4_lut (.A(databus_out[12]), .B(n10_c), .C(n2), .D(rw), .Z(databus[12])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfcfe;
    LUT4 i4_4_lut (.A(\read_value[12] ), .B(n8_c), .C(n1), .D(n28582), 
         .Z(n10_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut.init = 16'hfefc;
    LUT4 i2_4_lut (.A(\read_value[12]_adj_6 ), .B(read_value[12]), .C(n28451), 
         .D(n52), .Z(n8_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 n1016_bdd_3_lut_20539 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n27408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1016_bdd_3_lut_20539.init = 16'hcaca;
    LUT4 n1016_bdd_3_lut_20688 (.A(n1016), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n27409)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1016_bdd_3_lut_20688.init = 16'he2e2;
    LUT4 n986_bdd_3_lut_20655 (.A(n986), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n27464)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n986_bdd_3_lut_20655.init = 16'he2e2;
    LUT4 \register_1[[4__bdd_3_lut_20813  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n27994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_20813 .init = 16'hcaca;
    LUT4 register_addr_1__bdd_3_lut_20788 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n27992)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_20788.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_20787 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n27991)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_20787.init = 16'h2222;
    LUT4 \register_1[[4__bdd_2_lut_20814  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n27995)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_20814 .init = 16'h8888;
    LUT4 i5_4_lut_adj_70 (.A(databus_out[13]), .B(n10_adj_59), .C(n2_adj_8), 
         .D(rw), .Z(databus[13])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_70.init = 16'hfcfe;
    LUT4 i5_4_lut_adj_71 (.A(databus_out[9]), .B(n10_adj_61), .C(n2_adj_9), 
         .D(rw), .Z(databus[9])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_71.init = 16'hfcfe;
    LUT4 i5_4_lut_adj_72 (.A(databus_out[8]), .B(n10_adj_63), .C(n2_adj_10), 
         .D(rw), .Z(databus[8])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_72.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_73 (.A(\read_value[8]_adj_11 ), .B(n8_adj_65), .C(n1_adj_12), 
         .D(n28582), .Z(n10_adj_63)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_73.init = 16'hfefc;
    LUT4 i2_4_lut_adj_74 (.A(\read_value[8]_adj_13 ), .B(read_value[8]), 
         .C(n28451), .D(n52), .Z(n8_adj_65)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_74.init = 16'heca0;
    LUT4 i4_4_lut_adj_75 (.A(\read_value[9]_adj_14 ), .B(n8_adj_69), .C(n1_adj_15), 
         .D(n28582), .Z(n10_adj_61)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_75.init = 16'hfefc;
    LUT4 i2_4_lut_adj_76 (.A(read_size[0]), .B(\read_size[0]_adj_16 ), .C(\select[1] ), 
         .D(n28487), .Z(n9)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_76.init = 16'heca0;
    LUT4 i3_4_lut (.A(\read_size[0]_adj_17 ), .B(n28452), .C(n28476), 
         .D(\read_size[0]_adj_18 ), .Z(n10)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 i1_4_lut (.A(read_size_c[0]), .B(\read_size[0]_adj_19 ), .C(\select[7] ), 
         .D(\select[2] ), .Z(n8)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i4_4_lut_adj_77 (.A(n7), .B(\read_size[2]_adj_20 ), .C(n6_c), 
         .D(n28487), .Z(\reg_size[2] )) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_77.init = 16'hfefa;
    LUT4 i2_4_lut_adj_78 (.A(\read_size[2]_adj_21 ), .B(read_size[2]), .C(n28476), 
         .D(\select[1] ), .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_78.init = 16'heca0;
    LUT4 i1_4_lut_adj_79 (.A(\read_size[2]_adj_22 ), .B(\read_size[2]_adj_23 ), 
         .C(n28480), .D(n28452), .Z(n6_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_79.init = 16'heca0;
    LUT4 i14_2_lut_rep_447 (.A(\select[7] ), .B(rw), .Z(n28568)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam i14_2_lut_rep_447.init = 16'h8888;
    LUT4 Select_3961_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_292[0]), 
         .Z(n7_adj_82)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam Select_3961_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3958_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_292[3]), 
         .Z(n7_adj_83)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam Select_3958_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3959_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_292[2]), 
         .Z(n7_adj_84)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam Select_3959_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3957_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_292[4]), 
         .Z(n7_adj_85)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam Select_3957_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3956_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_292[5]), 
         .Z(n7_adj_86)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam Select_3956_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3955_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_292[6]), 
         .Z(n7_adj_87)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam Select_3955_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3954_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_292[7]), 
         .Z(n7_adj_88)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam Select_3954_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 n1001_bdd_3_lut_20665 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n27810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1001_bdd_3_lut_20665.init = 16'hcaca;
    LUT4 i7_4_lut (.A(n13), .B(n4), .C(n12), .D(n6_adj_89), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut_adj_80 (.A(\read_value[0]_adj_24 ), .B(n10_adj_91), .C(n7_adj_82), 
         .D(n28448), .Z(n13)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_80.init = 16'hfefc;
    LUT4 i4_4_lut_adj_81 (.A(\read_value[0]_adj_25 ), .B(\read_value[0]_adj_26 ), 
         .C(n28458), .D(n28582), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_81.init = 16'heca0;
    LUT4 Select_3961_i6_2_lut (.A(databus_out[0]), .B(rw), .Z(n6_adj_89)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3961_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_82 (.A(read_value[0]), .B(read_value_adj_146[0]), 
         .C(n52), .D(n64), .Z(n10_adj_91)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_82.init = 16'heca0;
    LUT4 i5_4_lut_adj_83 (.A(databus_out[31]), .B(n10_adj_96), .C(n2_adj_35), 
         .D(rw), .Z(databus[31])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_83.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_84 (.A(\read_value[9]_adj_36 ), .B(read_value[9]), 
         .C(n28451), .D(n52), .Z(n8_adj_69)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_84.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_20841 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n28233)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_20841.init = 16'he4e4;
    LUT4 i5_4_lut_adj_85 (.A(databus_out[21]), .B(n10_adj_100), .C(n2_adj_37), 
         .D(rw), .Z(databus[21])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_85.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_86 (.A(\read_value[21]_adj_38 ), .B(n8_adj_102), .C(n1_adj_39), 
         .D(n28582), .Z(n10_adj_100)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_86.init = 16'hfefc;
    LUT4 i4_4_lut_adj_87 (.A(\read_value[31]_adj_40 ), .B(n8_adj_104), .C(n1_adj_41), 
         .D(n28582), .Z(n10_adj_96)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_87.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_20840 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n28232)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_20840.init = 16'h2222;
    LUT4 \register_1[[5__bdd_3_lut_21386  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n28235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_21386 .init = 16'hcaca;
    LUT4 i2_4_lut_adj_88 (.A(\read_value[31]_adj_42 ), .B(read_value[31]), 
         .C(n28451), .D(n52), .Z(n8_adj_104)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_88.init = 16'heca0;
    LUT4 \register_1[[5__bdd_2_lut_21387  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n28236)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_21387 .init = 16'h8888;
    LUT4 i7_4_lut_adj_89 (.A(n13_adj_108), .B(n4_adj_43), .C(n12_adj_110), 
         .D(n6_adj_111), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_89.init = 16'hfffe;
    L6MUX21 i20563 (.D0(n27465), .D1(n27462), .SD(\register_addr[2] ), 
            .Z(n27466));
    LUT4 i5_4_lut_adj_90 (.A(\read_value[7]_adj_44 ), .B(n10_adj_113), .C(n7_adj_88), 
         .D(n28448), .Z(n13_adj_108)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_90.init = 16'hfefc;
    LUT4 Select_3969_i1_2_lut_rep_455 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n28576)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3969_i1_2_lut_rep_455.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n11943)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    FD1S3IX read_value__i7 (.D(n27829), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(n28387), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n28238), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n27997), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n27411), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n27813), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i2.GSR = "ENABLED";
    LUT4 i4_4_lut_adj_91 (.A(\read_value[13]_adj_45 ), .B(n8_adj_114), .C(n1_adj_46), 
         .D(n28582), .Z(n10_adj_59)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_91.init = 16'hfefc;
    FD1S3IX read_value__i1 (.D(n27466), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i7_4_lut_adj_92 (.A(n13_adj_116), .B(n4_adj_47), .C(n12_adj_118), 
         .D(n6_adj_119), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_92.init = 16'hfffe;
    LUT4 i5_4_lut_adj_93 (.A(\read_value[6]_adj_48 ), .B(n10_adj_121), .C(n7_adj_87), 
         .D(n28448), .Z(n13_adj_116)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_93.init = 16'hfefc;
    LUT4 i4_4_lut_adj_94 (.A(\read_value[7]_adj_49 ), .B(\read_value[7]_adj_50 ), 
         .C(n28458), .D(n28582), .Z(n12_adj_110)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_94.init = 16'heca0;
    LUT4 i2_4_lut_adj_95 (.A(\read_value[13]_adj_51 ), .B(read_value[13]), 
         .C(n28451), .D(n52), .Z(n8_adj_114)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_95.init = 16'heca0;
    LUT4 i4_4_lut_adj_96 (.A(\read_value[6]_adj_52 ), .B(\read_value[6]_adj_53 ), 
         .C(n28458), .D(n28582), .Z(n12_adj_118)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_96.init = 16'heca0;
    LUT4 Select_3955_i6_2_lut (.A(databus_out[6]), .B(rw), .Z(n6_adj_119)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3955_i6_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_97 (.A(databus_out[11]), .B(n10_adj_128), .C(n2_adj_54), 
         .D(rw), .Z(databus[11])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_97.init = 16'hfcfe;
    LUT4 Select_3954_i6_2_lut (.A(databus_out[7]), .B(rw), .Z(n6_adj_111)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3954_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_98 (.A(read_value[7]), .B(read_value_adj_146[7]), 
         .C(n52), .D(n64), .Z(n10_adj_113)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_98.init = 16'heca0;
    LUT4 i2_4_lut_adj_99 (.A(read_value[6]), .B(read_value_adj_146[6]), 
         .C(n52), .D(n64), .Z(n10_adj_121)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_99.init = 16'heca0;
    LUT4 i2_4_lut_adj_100 (.A(\read_value[21]_adj_55 ), .B(read_value[21]), 
         .C(n28451), .D(n52), .Z(n8_adj_102)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_100.init = 16'heca0;
    LUT4 n986_bdd_3_lut_20560 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n27463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n986_bdd_3_lut_20560.init = 16'hcaca;
    LUT4 register_addr_1__bdd_3_lut_20660 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n27689)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_20660.init = 16'he4e4;
    LUT4 i4_4_lut_adj_101 (.A(\read_value[11]_adj_56 ), .B(n8_adj_136), 
         .C(n1_adj_57), .D(n28582), .Z(n10_adj_128)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_101.init = 16'hfefc;
    LUT4 i2_4_lut_adj_102 (.A(\read_value[10]_adj_58 ), .B(read_value[10]), 
         .C(n28451), .D(n52), .Z(n8_adj_139)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_102.init = 16'heca0;
    PFUMX i20558 (.BLUT(n27461), .ALUT(n27460), .C0(\register_addr[1] ), 
          .Z(n27462));
    LUT4 n1001_bdd_3_lut_21090 (.A(n1001), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n27811)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1001_bdd_3_lut_21090.init = 16'he2e2;
    LUT4 i5_4_lut_adj_103 (.A(databus_out[30]), .B(n10_adj_140), .C(n2_adj_59), 
         .D(rw), .Z(databus[30])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_103.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_104 (.A(\read_value[30]_adj_60 ), .B(n8_adj_142), 
         .C(n1_adj_61), .D(n28582), .Z(n10_adj_140)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_104.init = 16'hfefc;
    LUT4 i7_4_lut_adj_105 (.A(n13_adj_144), .B(n4_adj_62), .C(n12_adj_146), 
         .D(n6_adj_147), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_105.init = 16'hfffe;
    LUT4 i5_4_lut_adj_106 (.A(\read_value[5]_adj_63 ), .B(n10_adj_149), 
         .C(n7_adj_86), .D(n28448), .Z(n13_adj_144)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_106.init = 16'hfefc;
    LUT4 i4_4_lut_adj_107 (.A(\read_value[5]_adj_64 ), .B(\read_value[5]_adj_65 ), 
         .C(n28458), .D(n28582), .Z(n12_adj_146)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_107.init = 16'heca0;
    LUT4 Select_3956_i6_2_lut (.A(databus_out[5]), .B(n30468), .Z(n6_adj_147)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3956_i6_2_lut.init = 16'h2222;
    L6MUX21 i20542 (.D0(n27410), .D1(n27407), .SD(\register_addr[2] ), 
            .Z(n27411));
    LUT4 i2_4_lut_adj_108 (.A(read_value[5]), .B(read_value_adj_146[5]), 
         .C(n52), .D(n64), .Z(n10_adj_149)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_108.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_20605 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n27460)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_20605.init = 16'h2222;
    LUT4 i2_4_lut_adj_109 (.A(\read_value[30]_adj_66 ), .B(read_value[30]), 
         .C(n28451), .D(n52), .Z(n8_adj_142)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_109.init = 16'heca0;
    LUT4 i7_4_lut_adj_110 (.A(n13_adj_156), .B(n4_adj_67), .C(n12_adj_158), 
         .D(n6_adj_159), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_110.init = 16'hfffe;
    LUT4 i5_4_lut_adj_111 (.A(\read_value[4]_adj_68 ), .B(n10_adj_161), 
         .C(n7_adj_85), .D(n28448), .Z(n13_adj_156)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_111.init = 16'hfefc;
    LUT4 i4_4_lut_adj_112 (.A(\read_value[4]_adj_69 ), .B(\read_value[4]_adj_70 ), 
         .C(n28458), .D(n28582), .Z(n12_adj_158)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_112.init = 16'heca0;
    L6MUX21 i20617 (.D0(n27693), .D1(n27690), .SD(\register_addr[2] ), 
            .Z(n27694));
    LUT4 Select_3957_i6_2_lut (.A(databus_out[4]), .B(rw), .Z(n6_adj_159)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3957_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_113 (.A(read_value[4]), .B(read_value_adj_146[4]), 
         .C(n52), .D(n64), .Z(n10_adj_161)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_113.init = 16'heca0;
    LUT4 i7_4_lut_adj_114 (.A(n13_adj_166), .B(n4_adj_71), .C(n12_adj_168), 
         .D(n6_adj_169), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_114.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_20606 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n27461)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_20606.init = 16'he4e4;
    LUT4 i5_4_lut_adj_115 (.A(\read_value[2]_adj_72 ), .B(n10_adj_171), 
         .C(n7_adj_84), .D(n28448), .Z(n13_adj_166)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_115.init = 16'hfefc;
    LUT4 i4_4_lut_adj_116 (.A(\read_value[2]_adj_73 ), .B(\read_value[2]_adj_74 ), 
         .C(n28458), .D(n28582), .Z(n12_adj_168)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_116.init = 16'heca0;
    L6MUX21 i20868 (.D0(n28386), .D1(n28383), .SD(\register_addr[2] ), 
            .Z(n28387));
    PFUMX i20866 (.BLUT(n28385), .ALUT(n28384), .C0(\register_addr[1] ), 
          .Z(n28386));
    PFUMX i20615 (.BLUT(n27692), .ALUT(n27691), .C0(\register_addr[1] ), 
          .Z(n27693));
    LUT4 Select_3959_i6_2_lut (.A(databus_out[2]), .B(rw), .Z(n6_adj_169)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3959_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_117 (.A(read_value[2]), .B(read_value_adj_146[2]), 
         .C(n52), .D(n64), .Z(n10_adj_171)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_117.init = 16'heca0;
    PFUMX i20863 (.BLUT(n28382), .ALUT(n28381), .C0(\register_addr[1] ), 
          .Z(n28383));
    PFUMX i20612 (.BLUT(n27689), .ALUT(n27688), .C0(\register_addr[1] ), 
          .Z(n27690));
    LUT4 i2_4_lut_adj_118 (.A(\read_value[11]_adj_75 ), .B(read_value[11]), 
         .C(n28451), .D(n52), .Z(n8_adj_136)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_118.init = 16'heca0;
    LUT4 n1046_bdd_3_lut_20985 (.A(n1046), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n27827)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1046_bdd_3_lut_20985.init = 16'he2e2;
    LUT4 i5_4_lut_adj_119 (.A(databus_out[28]), .B(n10_adj_178), .C(n2_adj_76), 
         .D(rw), .Z(databus[28])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_119.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_120 (.A(\read_value[28]_adj_77 ), .B(n8_adj_180), 
         .C(n1_adj_78), .D(n28582), .Z(n10_adj_178)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_120.init = 16'hfefc;
    LUT4 i2_4_lut_adj_121 (.A(\read_value[28]_adj_79 ), .B(read_value[28]), 
         .C(n28451), .D(n52), .Z(n8_adj_180)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_121.init = 16'heca0;
    LUT4 i5_4_lut_adj_122 (.A(databus_out[27]), .B(n10_adj_184), .C(n2_adj_80), 
         .D(rw), .Z(databus[27])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_122.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_123 (.A(\read_value[27]_adj_81 ), .B(n8_adj_186), 
         .C(n1_adj_82), .D(n28582), .Z(n10_adj_184)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_123.init = 16'hfefc;
    LUT4 i7_4_lut_adj_124 (.A(n1_adj_83), .B(n14), .C(n10_adj_189), .D(n7_adj_190), 
         .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_124.init = 16'hfffe;
    LUT4 i5_4_lut_adj_125 (.A(databus_out[10]), .B(n10_adj_191), .C(n2_adj_84), 
         .D(rw), .Z(databus[10])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_125.init = 16'hfcfe;
    LUT4 i6_4_lut (.A(\read_value[1]_adj_85 ), .B(n12_adj_194), .C(n6), 
         .D(n28451), .Z(n14)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 i5_4_lut_adj_126 (.A(databus_out[20]), .B(n10_adj_196), .C(n2_adj_86), 
         .D(rw), .Z(databus[20])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_126.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_127 (.A(\read_value[20]_adj_87 ), .B(n8_adj_198), 
         .C(n1_adj_88), .D(n28582), .Z(n10_adj_196)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_127.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_20671 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n27807)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_20671.init = 16'h2222;
    LUT4 i2_4_lut_adj_128 (.A(\read_value[27]_adj_89 ), .B(read_value[27]), 
         .C(n28451), .D(n52), .Z(n8_adj_186)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_128.init = 16'heca0;
    LUT4 i5_4_lut_adj_129 (.A(databus_out[14]), .B(n10_adj_202), .C(n2_adj_90), 
         .D(rw), .Z(databus[14])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_129.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_130 (.A(\read_value[20]_adj_91 ), .B(read_value[20]), 
         .C(n28451), .D(n52), .Z(n8_adj_198)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_130.init = 16'heca0;
    LUT4 i5_4_lut_adj_131 (.A(databus_out[19]), .B(n10_adj_206), .C(n2_adj_92), 
         .D(rw), .Z(databus[19])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_131.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_132 (.A(\read_value[14]_adj_93 ), .B(n8_adj_208), 
         .C(n1_adj_94), .D(n28582), .Z(n10_adj_202)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_132.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_20672 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n27808)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_20672.init = 16'he4e4;
    LUT4 i2_4_lut_adj_133 (.A(\read_value[14]_adj_95 ), .B(read_value[14]), 
         .C(n28451), .D(n52), .Z(n8_adj_208)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_133.init = 16'heca0;
    LUT4 i2_4_lut_adj_134 (.A(read_value[1]), .B(read_value_adj_146[1]), 
         .C(n52), .D(n64), .Z(n10_adj_189)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_134.init = 16'heca0;
    L6MUX21 i20793 (.D0(n28237), .D1(n28234), .SD(\register_addr[2] ), 
            .Z(n28238));
    LUT4 i4_4_lut_adj_135 (.A(\read_value[19]_adj_96 ), .B(n8_adj_214), 
         .C(n1_adj_97), .D(n28582), .Z(n10_adj_206)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_135.init = 16'hfefc;
    PFUMX i20791 (.BLUT(n28236), .ALUT(n28235), .C0(\register_addr[1] ), 
          .Z(n28237));
    FD1S3IX read_value__i0 (.D(n27694), .CK(\select[7] ), .CD(n28439), 
            .Q(read_value_adj_292[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=621, LSE_RLINE=633 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i7_4_lut_adj_136 (.A(n13_adj_216), .B(n4_adj_98), .C(n12_adj_218), 
         .D(n6_adj_219), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_136.init = 16'hfffe;
    PFUMX i20789 (.BLUT(n28233), .ALUT(n28232), .C0(\register_addr[1] ), 
          .Z(n28234));
    LUT4 i4_4_lut_adj_137 (.A(\read_value[10]_adj_99 ), .B(n8_adj_139), 
         .C(n1_adj_100), .D(n28582), .Z(n10_adj_191)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_137.init = 16'hfefc;
    LUT4 Select_3960_i7_2_lut (.A(databus_out[1]), .B(n30468), .Z(n7_adj_190)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3960_i7_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_138 (.A(\read_value[3]_adj_101 ), .B(n10_adj_223), 
         .C(n7_adj_83), .D(n28448), .Z(n13_adj_216)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_138.init = 16'hfefc;
    LUT4 i5_4_lut_adj_139 (.A(databus_out[26]), .B(n10_adj_224), .C(n2_adj_102), 
         .D(rw), .Z(databus[26])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_139.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_140 (.A(\read_value[19]_adj_103 ), .B(read_value[19]), 
         .C(n28451), .D(n52), .Z(n8_adj_214)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_140.init = 16'heca0;
    LUT4 i4_4_lut_adj_141 (.A(\read_value[26]_adj_104 ), .B(n8_adj_228), 
         .C(n1_adj_105), .D(n28582), .Z(n10_adj_224)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_141.init = 16'hfefc;
    LUT4 i4_4_lut_adj_142 (.A(\read_value[3]_adj_106 ), .B(\read_value[3]_adj_107 ), 
         .C(n28458), .D(n28582), .Z(n12_adj_218)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_142.init = 16'heca0;
    LUT4 i2_4_lut_adj_143 (.A(\read_value[26]_adj_108 ), .B(read_value[26]), 
         .C(n28451), .D(n52), .Z(n8_adj_228)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_143.init = 16'heca0;
    LUT4 Select_3958_i6_2_lut (.A(databus_out[3]), .B(n30468), .Z(n6_adj_219)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3958_i6_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_144 (.A(databus_out[25]), .B(n10_adj_234), .C(n2_adj_109), 
         .D(rw), .Z(databus[25])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_144.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_145 (.A(\read_value[25]_adj_110 ), .B(n8_adj_236), 
         .C(n1_adj_111), .D(n28582), .Z(n10_adj_234)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_145.init = 16'hfefc;
    LUT4 i5_4_lut_adj_146 (.A(databus_out[18]), .B(n10_adj_238), .C(n2_adj_112), 
         .D(rw), .Z(databus[18])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_146.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_147 (.A(\read_value[18]_adj_113 ), .B(n8_adj_240), 
         .C(n1_adj_114), .D(n28582), .Z(n10_adj_238)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_147.init = 16'hfefc;
    LUT4 i2_4_lut_adj_148 (.A(\read_value[25]_adj_115 ), .B(read_value[25]), 
         .C(n28451), .D(n52), .Z(n8_adj_236)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_148.init = 16'heca0;
    LUT4 i2_4_lut_adj_149 (.A(\read_value[18]_adj_116 ), .B(read_value[18]), 
         .C(n28451), .D(n52), .Z(n8_adj_240)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_149.init = 16'heca0;
    LUT4 i2_4_lut_adj_150 (.A(read_value[3]), .B(read_value_adj_146[3]), 
         .C(n52), .D(n64), .Z(n10_adj_223)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_150.init = 16'heca0;
    LUT4 i5_4_lut_adj_151 (.A(databus_out[17]), .B(n10_adj_248), .C(n2_adj_117), 
         .D(rw), .Z(databus[17])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_151.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_152 (.A(\read_value[17]_adj_118 ), .B(n8_adj_250), 
         .C(n1_adj_119), .D(n28582), .Z(n10_adj_248)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_152.init = 16'hfefc;
    LUT4 i2_4_lut_adj_153 (.A(\read_value[17]_adj_120 ), .B(read_value[17]), 
         .C(n28451), .D(n52), .Z(n8_adj_250)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_153.init = 16'heca0;
    LUT4 i5_4_lut_adj_154 (.A(databus_out[24]), .B(n10_adj_254), .C(n2_adj_121), 
         .D(rw), .Z(databus[24])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_154.init = 16'hfcfe;
    L6MUX21 i20729 (.D0(n27996), .D1(n27993), .SD(\register_addr[2] ), 
            .Z(n27997));
    LUT4 i4_4_lut_adj_155 (.A(\read_value[24]_adj_122 ), .B(n8_adj_256), 
         .C(n1_adj_123), .D(n28582), .Z(n10_adj_254)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_155.init = 16'hfefc;
    PFUMX i20727 (.BLUT(n27995), .ALUT(n27994), .C0(\register_addr[1] ), 
          .Z(n27996));
    LUT4 i2_4_lut_adj_156 (.A(\read_value[24]_adj_124 ), .B(read_value[24]), 
         .C(n28451), .D(n52), .Z(n8_adj_256)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_156.init = 16'heca0;
    PFUMX i20540 (.BLUT(n27409), .ALUT(n27408), .C0(\register_addr[1] ), 
          .Z(n27410));
    LUT4 i4_4_lut_adj_157 (.A(\read_value[1]_adj_125 ), .B(read_value_adj_292[1]), 
         .C(n28458), .D(n28568), .Z(n12_adj_194)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_157.init = 16'heca0;
    LUT4 i5_4_lut_adj_158 (.A(databus_out[16]), .B(n10_adj_261), .C(n2_adj_126), 
         .D(rw), .Z(databus[16])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_158.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_159 (.A(\read_value[16]_adj_127 ), .B(n8_adj_263), 
         .C(n1_adj_128), .D(n28582), .Z(n10_adj_261)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_159.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_20711 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n27823)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_20711.init = 16'h2222;
    LUT4 i5_4_lut_adj_160 (.A(databus_out[23]), .B(n10_adj_265), .C(n2_adj_129), 
         .D(rw), .Z(databus[23])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_160.init = 16'hfcfe;
    PFUMX i20725 (.BLUT(n27992), .ALUT(n27991), .C0(\register_addr[1] ), 
          .Z(n27993));
    LUT4 i5_4_lut_adj_161 (.A(databus_out[29]), .B(n10_adj_267), .C(n2_adj_130), 
         .D(rw), .Z(databus[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_161.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_162 (.A(\read_value[29]_adj_131 ), .B(n8_adj_269), 
         .C(n1_adj_132), .D(n28582), .Z(n10_adj_267)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_162.init = 16'hfefc;
    LUT4 i2_4_lut_adj_163 (.A(\read_value[16]_adj_133 ), .B(read_value[16]), 
         .C(n28451), .D(n52), .Z(n8_adj_263)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_163.init = 16'heca0;
    LUT4 i2_4_lut_adj_164 (.A(\read_value[29]_adj_134 ), .B(read_value[29]), 
         .C(n28451), .D(n52), .Z(n8_adj_269)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_164.init = 16'heca0;
    LUT4 i4_4_lut_adj_165 (.A(\read_value[23]_adj_135 ), .B(n8_adj_275), 
         .C(n1_adj_136), .D(n28582), .Z(n10_adj_265)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_165.init = 16'hfefc;
    LUT4 i5_4_lut_adj_166 (.A(databus_out[15]), .B(n10_adj_277), .C(n2_adj_137), 
         .D(rw), .Z(databus[15])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_166.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_167 (.A(\read_value[23]_adj_138 ), .B(read_value[23]), 
         .C(n28451), .D(n52), .Z(n8_adj_275)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_167.init = 16'heca0;
    LUT4 i4_4_lut_adj_168 (.A(\read_value[15]_adj_139 ), .B(n8_adj_281), 
         .C(n1_adj_140), .D(n28582), .Z(n10_adj_277)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_168.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_20712 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n27824)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_20712.init = 16'he4e4;
    LUT4 i5_4_lut_adj_169 (.A(databus_out[22]), .B(n10_adj_283), .C(n2_adj_141), 
         .D(rw), .Z(databus[22])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_169.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_170 (.A(\read_value[22]_adj_142 ), .B(n8_adj_285), 
         .C(n1_adj_143), .D(n28582), .Z(n10_adj_283)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_170.init = 16'hfefc;
    LUT4 i2_4_lut_adj_171 (.A(\read_value[15]_adj_144 ), .B(read_value[15]), 
         .C(n28451), .D(n52), .Z(n8_adj_281)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_171.init = 16'heca0;
    PFUMX i20537 (.BLUT(n27406), .ALUT(n27405), .C0(\register_addr[1] ), 
          .Z(n27407));
    LUT4 i2_4_lut_adj_172 (.A(\read_value[22]_adj_145 ), .B(read_value[22]), 
         .C(n28451), .D(n52), .Z(n8_adj_285)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_172.init = 16'heca0;
    PFUMX i20561 (.BLUT(n27464), .ALUT(n27463), .C0(\register_addr[1] ), 
          .Z(n27465));
    PWMReceiver recv_ch8 (.debug_c_c(debug_c_c), .n30470(n30470), .rc_ch8_c(rc_ch8_c), 
            .GND_net(GND_net), .n26922(n26922), .n30469(n30469), .n26942(n26942), 
            .\register[6] ({\register[6] }), .n12605(n12605), .n1046(n1046), 
            .n24743(n24743)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(257[14] 261[36])
    PWMReceiver_U1 recv_ch7 (.GND_net(GND_net), .debug_c_c(debug_c_c), .n30471(n30471), 
            .n30470(n30470), .\register[5] ({\register[5] }), .n13489(n13489), 
            .rc_ch7_c(rc_ch7_c), .n26949(n26949), .n1031(n1031), .n24707(n24707), 
            .n27040(n27040), .n30469(n30469)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(252[14] 256[36])
    PWMReceiver_U2 recv_ch4 (.debug_c_c(debug_c_c), .n30471(n30471), .GND_net(GND_net), 
            .\register[4] ({\register[4] }), .n13527(n13527), .n30470(n30470), 
            .rc_ch4_c(rc_ch4_c), .n26947(n26947), .n1016(n1016), .n24721(n24721), 
            .n27035(n27035), .n30469(n30469)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(247[14] 251[36])
    PWMReceiver_U3 recv_ch3 (.debug_c_c(debug_c_c), .n30471(n30471), .GND_net(GND_net), 
            .\register[3] ({\register[3] }), .n13534(n13534), .n30470(n30470), 
            .rc_ch3_c(rc_ch3_c), .n27027(n27027), .n30469(n30469), .n26939(n26939), 
            .n1001(n1001), .n24755(n24755)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(242[14] 246[36])
    PWMReceiver_U4 recv_ch2 (.GND_net(GND_net), .debug_c_c(debug_c_c), .n30470(n30470), 
            .rc_ch2_c(rc_ch2_c), .n26945(n26945), .\register[2] ({\register[2] }), 
            .n13535(n13535), .n986(n986), .n24741(n24741), .n27025(n27025), 
            .n30469(n30469), .n28403(n28403), .n30471(n30471)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(237[14] 241[36])
    PWMReceiver_U5 recv_ch1 (.debug_c_c(debug_c_c), .n30470(n30470), .n26907(n26907), 
            .rc_ch1_c(rc_ch1_c), .GND_net(GND_net), .\register[1] ({\register[1] }), 
            .n13536(n13536), .n971(n971), .n24716(n24716), .n27023(n27023), 
            .n30469(n30469)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(232[17] 236[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (debug_c_c, n30470, rc_ch8_c, GND_net, n26922, 
            n30469, n26942, \register[6] , n12605, n1046, n24743) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30470;
    input rc_ch8_c;
    input GND_net;
    output n26922;
    input n30469;
    output n26942;
    output [7:0]\register[6] ;
    input n12605;
    output n1046;
    input n24743;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n28488, n28516, n28454, n26292;
    wire [7:0]n944;
    wire [7:0]n43;
    
    wire n28522, n6, n4, n28523, n5, n24923, n26621, n28515, 
        n1052, n1040, n28416, n30465, n26620, n26548, n28453, 
        n28483, n28427, n28426, n26622, n10, n24064, n16, n14707, 
        n26, n24063, n28521, n11696, n8, n33, n28484, n4_adj_54, 
        n28456, n24062, n24061, n5_adj_55, n26721, n23868;
    wire [15:0]n116;
    
    wire n23867, n23866, n23865, n23864, n24742, n23863, n23862, 
        n23861, n4_adj_56;
    
    LUT4 i1_2_lut_rep_367_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n28488)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_367_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_333_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n28516), 
         .D(count[0]), .Z(n28454)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_333_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(n26292), .B(n944[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i2687_2_lut_rep_401 (.A(count[1]), .B(count[2]), .Z(n28522)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2687_2_lut_rep_401.init = 16'h8888;
    LUT4 i4_3_lut_rep_395_4_lut (.A(count[1]), .B(count[2]), .C(n6), .D(count[3]), 
         .Z(n28516)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_3_lut_rep_395_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_402 (.A(count[15]), .B(count[14]), .Z(n28523)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_402.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n24923), 
         .Z(n26621)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i19970_2_lut_rep_394_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n28515)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i19970_2_lut_rep_394_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_58 (.A(n26292), .B(n944[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_58.init = 16'h4444;
    LUT4 i1_2_lut_adj_59 (.A(n26292), .B(n944[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_59.init = 16'h4444;
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n30470), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1052));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1052), .SP(n30470), .CK(debug_c_c), .Q(n1040));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i20304_3_lut_3_lut_4_lut (.A(n28523), .B(n24923), .C(n28416), 
         .D(n30465), .Z(n26620)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i20304_3_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_60 (.A(n26292), .B(n944[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_60.init = 16'h4444;
    LUT4 i1_2_lut_rep_332_4_lut (.A(n28515), .B(count[13]), .C(n26548), 
         .D(count[9]), .Z(n28453)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_332_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_306_3_lut (.A(count[9]), .B(n28483), .C(count[8]), 
         .Z(n28427)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_306_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_61 (.A(n26292), .B(n944[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_61.init = 16'h4444;
    LUT4 i20323_4_lut (.A(n28426), .B(n26622), .C(n26292), .D(n10), 
         .Z(n26922)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i20323_4_lut.init = 16'h3323;
    CCU2D sub_59_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24064), 
          .S0(n944[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_59_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_9.INIT1 = 16'h0000;
    defparam sub_59_add_2_9.INJECT1_0 = "NO";
    defparam sub_59_add_2_9.INJECT1_1 = "NO";
    LUT4 i8_4_lut (.A(n28515), .B(n16), .C(count[13]), .D(count[11]), 
         .Z(n14707)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i8_4_lut.init = 16'h0004;
    LUT4 i7_4_lut (.A(count[10]), .B(n30469), .C(n26), .D(n26622), .Z(n16)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i7_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_adj_62 (.A(n26292), .B(n944[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_62.init = 16'h4444;
    CCU2D sub_59_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24063), 
          .COUT(n24064), .S0(n944[5]), .S1(n944[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_59_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_7.INJECT1_0 = "NO";
    defparam sub_59_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n28453), .B(count[8]), .C(n28521), .D(n28516), 
         .Z(n26292)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfbbb;
    LUT4 i13290_4_lut (.A(n11696), .B(count[1]), .C(n6), .D(n8), .Z(n33)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i13290_4_lut.init = 16'hfaea;
    LUT4 i3_3_lut (.A(count[2]), .B(count[3]), .C(count[0]), .Z(n8)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut (.A(count[7]), .B(count[8]), .C(count[6]), .Z(n11696)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_63 (.A(count[5]), .B(count[4]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_adj_63.init = 16'h8888;
    LUT4 i10_3_lut_4_lut_4_lut (.A(n28484), .B(n28521), .C(n4_adj_54), 
         .D(n28427), .Z(n10)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i10_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_adj_64 (.A(n1052), .B(n1040), .Z(n26622)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_64.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_65 (.A(count[4]), .B(count[5]), .C(count[3]), .D(n28522), 
         .Z(n4_adj_54)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_65.init = 16'hccc8;
    LUT4 i1_2_lut_rep_335_3_lut_4_lut (.A(count[8]), .B(n28521), .C(n28516), 
         .D(count[0]), .Z(n28456)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_335_3_lut_4_lut.init = 16'h8000;
    LUT4 i33_3_lut_4_lut (.A(n28484), .B(n28488), .C(count[9]), .D(n33), 
         .Z(n26)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_3_lut_4_lut.init = 16'h08f8;
    CCU2D sub_59_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24062), 
          .COUT(n24063), .S0(n944[3]), .S1(n944[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_59_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_5.INJECT1_0 = "NO";
    defparam sub_59_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24061), 
          .COUT(n24062), .S0(n944[1]), .S1(n944[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_59_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_3.INJECT1_0 = "NO";
    defparam sub_59_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24061), 
          .S1(n944[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_59_add_2_1.INIT0 = 16'hF000;
    defparam sub_59_add_2_1.INIT1 = 16'h5555;
    defparam sub_59_add_2_1.INJECT1_0 = "NO";
    defparam sub_59_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_66 (.A(n26292), .B(n944[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_66.init = 16'h4444;
    LUT4 i13683_2_lut (.A(n944[7]), .B(n26292), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13683_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_4_lut (.A(n28456), .B(n30465), .C(n28453), .D(n26292), 
         .Z(n5_adj_55)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    LUT4 i1_3_lut_rep_295_4_lut (.A(count[8]), .B(n28453), .C(n4_adj_54), 
         .D(n28521), .Z(n28416)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_3_lut_rep_295_4_lut.init = 16'hfeee;
    LUT4 i20031_3_lut_4_lut (.A(count[8]), .B(n28453), .C(n4_adj_54), 
         .D(n28454), .Z(n26721)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i20031_3_lut_4_lut.init = 16'hfeee;
    CCU2D add_1618_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n23868), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_17.INIT0 = 16'hd222;
    defparam add_1618_17.INIT1 = 16'h0000;
    defparam add_1618_17.INJECT1_0 = "NO";
    defparam add_1618_17.INJECT1_1 = "NO";
    CCU2D add_1618_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23867), 
          .COUT(n23868), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_15.INIT0 = 16'hd222;
    defparam add_1618_15.INIT1 = 16'hd222;
    defparam add_1618_15.INJECT1_0 = "NO";
    defparam add_1618_15.INJECT1_1 = "NO";
    CCU2D add_1618_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23866), 
          .COUT(n23867), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_13.INIT0 = 16'hd222;
    defparam add_1618_13.INIT1 = 16'hd222;
    defparam add_1618_13.INJECT1_0 = "NO";
    defparam add_1618_13.INJECT1_1 = "NO";
    CCU2D add_1618_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23865), 
          .COUT(n23866), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_11.INIT0 = 16'hd222;
    defparam add_1618_11.INIT1 = 16'hd222;
    defparam add_1618_11.INJECT1_0 = "NO";
    defparam add_1618_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_67 (.A(count[11]), .B(count[10]), .Z(n26548)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_67.init = 16'heeee;
    LUT4 i21_3_lut_rep_305_4_lut_4_lut (.A(count[9]), .B(n28483), .C(n33), 
         .D(n28456), .Z(n28426)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(D)))) */ ;
    defparam i21_3_lut_rep_305_4_lut_4_lut.init = 16'h1302;
    LUT4 i13765_3_lut_rep_462 (.A(count[9]), .B(n28483), .C(n33), .Z(n30465)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i13765_3_lut_rep_462.init = 16'hecec;
    CCU2D add_1618_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23864), 
          .COUT(n23865), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_9.INIT0 = 16'hd222;
    defparam add_1618_9.INIT1 = 16'hd222;
    defparam add_1618_9.INJECT1_0 = "NO";
    defparam add_1618_9.INJECT1_1 = "NO";
    LUT4 i3_3_lut_rep_362_4_lut (.A(count[12]), .B(n28523), .C(n26548), 
         .D(count[13]), .Z(n28483)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_362_4_lut.init = 16'hfffe;
    LUT4 i20343_4_lut (.A(n28523), .B(n5), .C(n24923), .D(n24742), .Z(n26942)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i20343_4_lut.init = 16'h3233;
    LUT4 i1_2_lut_rep_363_4_lut (.A(n28522), .B(count[3]), .C(n6), .D(count[0]), 
         .Z(n28484)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_363_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_68 (.A(n5_adj_55), .B(n26622), .C(n26721), .D(n30465), 
         .Z(n24742)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_68.init = 16'hccec;
    CCU2D add_1618_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23863), 
          .COUT(n23864), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_7.INIT0 = 16'hd222;
    defparam add_1618_7.INIT1 = 16'hd222;
    defparam add_1618_7.INJECT1_0 = "NO";
    defparam add_1618_7.INJECT1_1 = "NO";
    CCU2D add_1618_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23862), 
          .COUT(n23863), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_5.INIT0 = 16'hd222;
    defparam add_1618_5.INIT1 = 16'hd222;
    defparam add_1618_5.INJECT1_0 = "NO";
    defparam add_1618_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_400 (.A(count[7]), .B(count[6]), .Z(n28521)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_400.init = 16'h8888;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    CCU2D add_1618_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23861), 
          .COUT(n23862), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_3.INIT0 = 16'hd222;
    defparam add_1618_3.INIT1 = 16'hd222;
    defparam add_1618_3.INJECT1_0 = "NO";
    defparam add_1618_3.INJECT1_1 = "NO";
    CCU2D add_1618_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n26621), .B1(n1052), .C1(count[0]), .D1(n1040), .COUT(n23861), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1618_1.INIT0 = 16'hF000;
    defparam add_1618_1.INIT1 = 16'ha565;
    defparam add_1618_1.INJECT1_0 = "NO";
    defparam add_1618_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3AX valid_48 (.D(n26620), .SP(n24743), .CK(debug_c_c), .Q(n1046));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12605), .PD(n14707), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(n1040), .B(n1052), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n26548), .D(n4_adj_56), 
         .Z(n24923)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_69 (.A(count[5]), .B(count[9]), .C(n28488), .D(n4), 
         .Z(n4_adj_56)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_69.init = 16'hfcec;
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (GND_net, debug_c_c, n30471, n30470, \register[5] , 
            n13489, rc_ch7_c, n26949, n1031, n24707, n27040, n30469) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n30471;
    input n30470;
    output [7:0]\register[5] ;
    input n13489;
    input rc_ch7_c;
    output n26949;
    output n1031;
    input n24707;
    output n27040;
    input n30469;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n28524, n5, n24924, n26602, n28525, n28490, n5_adj_49, 
        n111, n103, n28526, n28460, n4, n28527, n6, n28489, 
        n28528, n26780, n28461, n4_adj_50, n28417, n23875;
    wire [15:0]n116;
    
    wire n23876, n23874, n23873, n12439, n154, n26740, n14918;
    wire [7:0]n43;
    
    wire n23872, n23871, n1037;
    wire [7:0]n935;
    
    wire n26294, n24068, n24067, n24066, n24065, n28433, n28432, 
        n26735, n10, n23870, n26603, n23869, n1025, n152, n24706, 
        n5_adj_51, n26708, n54, n4_adj_52, n6_adj_53, n26484, n11;
    
    LUT4 i1_2_lut_rep_403 (.A(count[15]), .B(count[14]), .Z(n28524)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_403.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n24924), 
         .Z(n26602)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_404 (.A(count[4]), .B(count[5]), .Z(n28525)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_404.init = 16'h8888;
    LUT4 i1_2_lut_rep_369_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n28490)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_369_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n5_adj_49)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[4]), .B(count[5]), .C(n111), .Z(n103)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i2_2_lut_rep_339_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(n28526), 
         .D(count[3]), .Z(n28460)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut_rep_339_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_405 (.A(count[2]), .B(count[1]), .Z(n28526)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_405.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(n28527), 
         .D(count[8]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_406 (.A(count[7]), .B(count[6]), .Z(n28527)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_406.init = 16'h8888;
    LUT4 i1_2_lut_rep_368_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n28489)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_368_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_407 (.A(count[11]), .B(count[10]), .Z(n28528)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_407.init = 16'heeee;
    LUT4 i20086_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n26780)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20086_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_rep_296_4_lut (.A(count[8]), .B(n28461), .C(n4_adj_50), 
         .D(n28527), .Z(n28417)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_3_lut_rep_296_4_lut.init = 16'hfeee;
    CCU2D add_1614_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23875), 
          .COUT(n23876), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_15.INIT0 = 16'hd222;
    defparam add_1614_15.INIT1 = 16'hd222;
    defparam add_1614_15.INJECT1_0 = "NO";
    defparam add_1614_15.INJECT1_1 = "NO";
    CCU2D add_1614_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23874), 
          .COUT(n23875), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_13.INIT0 = 16'hd222;
    defparam add_1614_13.INIT1 = 16'hd222;
    defparam add_1614_13.INJECT1_0 = "NO";
    defparam add_1614_13.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    CCU2D add_1614_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23873), 
          .COUT(n23874), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_11.INIT0 = 16'hd222;
    defparam add_1614_11.INIT1 = 16'hd222;
    defparam add_1614_11.INJECT1_0 = "NO";
    defparam add_1614_11.INJECT1_1 = "NO";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    LUT4 i20046_3_lut (.A(n12439), .B(count[9]), .C(n154), .Z(n26740)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i20046_3_lut.init = 16'heaea;
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1614_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23872), 
          .COUT(n23873), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_9.INIT0 = 16'hd222;
    defparam add_1614_9.INIT1 = 16'hd222;
    defparam add_1614_9.INJECT1_0 = "NO";
    defparam add_1614_9.INJECT1_1 = "NO";
    CCU2D add_1614_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23871), 
          .COUT(n23872), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_7.INIT0 = 16'hd222;
    defparam add_1614_7.INIT1 = 16'hd222;
    defparam add_1614_7.INJECT1_0 = "NO";
    defparam add_1614_7.INJECT1_1 = "NO";
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n30470), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1037));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i13464_2_lut (.A(n935[0]), .B(n26294), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13464_2_lut.init = 16'h2222;
    CCU2D sub_58_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24068), 
          .S0(n935[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_58_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_9.INIT1 = 16'h0000;
    defparam sub_58_add_2_9.INJECT1_0 = "NO";
    defparam sub_58_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24067), 
          .COUT(n24068), .S0(n935[5]), .S1(n935[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_58_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_7.INJECT1_0 = "NO";
    defparam sub_58_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24066), 
          .COUT(n24067), .S0(n935[3]), .S1(n935[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_58_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_5.INJECT1_0 = "NO";
    defparam sub_58_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24065), 
          .COUT(n24066), .S0(n935[1]), .S1(n935[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_58_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_3.INJECT1_0 = "NO";
    defparam sub_58_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24065), 
          .S1(n935[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_58_add_2_1.INIT0 = 16'hF000;
    defparam sub_58_add_2_1.INIT1 = 16'h5555;
    defparam sub_58_add_2_1.INJECT1_0 = "NO";
    defparam sub_58_add_2_1.INJECT1_1 = "NO";
    LUT4 i20041_3_lut_4_lut (.A(n28527), .B(n28433), .C(n4_adj_50), .D(n28432), 
         .Z(n26735)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i20041_3_lut_4_lut.init = 16'hff80;
    LUT4 i10_3_lut_4_lut_4_lut (.A(n28527), .B(n28432), .C(n4_adj_50), 
         .D(n28433), .Z(n10)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i10_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_312_3_lut_4_lut (.A(count[3]), .B(n28525), .C(count[0]), 
         .D(n28526), .Z(n28433)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_312_3_lut_4_lut.init = 16'h8000;
    CCU2D add_1614_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23870), 
          .COUT(n23871), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_5.INIT0 = 16'hd222;
    defparam add_1614_5.INIT1 = 16'hd222;
    defparam add_1614_5.INJECT1_0 = "NO";
    defparam add_1614_5.INJECT1_1 = "NO";
    LUT4 i20388_3_lut_3_lut_4_lut (.A(n28524), .B(n24924), .C(n28417), 
         .D(n26740), .Z(n26603)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i20388_3_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D add_1614_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n23869), 
          .COUT(n23870), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_3.INIT0 = 16'hd222;
    defparam add_1614_3.INIT1 = 16'hd222;
    defparam add_1614_3.INJECT1_0 = "NO";
    defparam add_1614_3.INJECT1_1 = "NO";
    CCU2D add_1614_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n26602), .B1(n1037), .C1(count[0]), .D1(n1025), .COUT(n23869), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_1.INIT0 = 16'hF000;
    defparam add_1614_1.INIT1 = 16'ha565;
    defparam add_1614_1.INJECT1_0 = "NO";
    defparam add_1614_1.INJECT1_1 = "NO";
    LUT4 i13681_2_lut (.A(n935[6]), .B(n26294), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13681_2_lut.init = 16'h2222;
    PFUMX i12474 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    LUT4 i5_2_lut (.A(n1025), .B(n1037), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i20350_4_lut (.A(n28524), .B(n5), .C(n24924), .D(n24706), .Z(n26949)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i20350_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5_adj_51), .B(n26708), .C(n26735), .D(n26740), 
         .Z(n24706)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i1_2_lut (.A(n54), .B(n26294), .Z(n5_adj_51)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    FD1P3AX prev_in_46 (.D(n1037), .SP(n30470), .CK(debug_c_c), .Q(n1025));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i13680_2_lut (.A(n935[5]), .B(n26294), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13680_2_lut.init = 16'h2222;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n28528), .D(n4_adj_52), 
         .Z(n24924)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_53 (.A(count[9]), .B(count[4]), .C(n28489), .D(n4), 
         .Z(n4_adj_52)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_53.init = 16'hfaea;
    LUT4 i23_4_lut (.A(n111), .B(count[2]), .C(n28525), .D(n6_adj_53), 
         .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6_adj_53)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n111)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_54 (.A(n28490), .B(n28526), .C(n28489), 
         .D(count[0]), .Z(n26484)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_54.init = 16'h8000;
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13489), .PD(n14918), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i13679_2_lut (.A(n935[4]), .B(n26294), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13679_2_lut.init = 16'h2222;
    LUT4 i13678_2_lut (.A(n935[3]), .B(n26294), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13678_2_lut.init = 16'h2222;
    FD1P3IX valid_48 (.D(n26603), .SP(n24707), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1031));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_340 (.A(count[9]), .B(n12439), .Z(n28461)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_340.init = 16'heeee;
    LUT4 i1_2_lut_rep_311_3_lut (.A(count[9]), .B(n12439), .C(count[8]), 
         .Z(n28432)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_311_3_lut.init = 16'hfefe;
    LUT4 i13677_2_lut (.A(n935[2]), .B(n26294), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13677_2_lut.init = 16'h2222;
    LUT4 i13676_2_lut (.A(n935[1]), .B(n26294), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13676_2_lut.init = 16'h2222;
    LUT4 i20441_4_lut (.A(n54), .B(n26708), .C(n26294), .D(n10), .Z(n27040)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i20441_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_55 (.A(n30469), .B(n28524), .C(n11), .D(n26780), 
         .Z(n14918)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_55.init = 16'h0020;
    LUT4 i4_4_lut (.A(n26484), .B(n26708), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i13682_2_lut (.A(n935[7]), .B(n26294), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i13682_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_56 (.A(n28461), .B(count[8]), .C(n28527), .D(n28460), 
         .Z(n26294)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_56.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n28524), .D(n28528), 
         .Z(n12439)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_57 (.A(count[5]), .B(count[3]), .C(count[4]), .D(n28526), 
         .Z(n4_adj_50)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_57.init = 16'haaa8;
    LUT4 i21_4_lut (.A(n5_adj_49), .B(n26740), .C(n28461), .D(n6), .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    CCU2D add_1614_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n23876), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1614_17.INIT0 = 16'hd222;
    defparam add_1614_17.INIT1 = 16'h0000;
    defparam add_1614_17.INJECT1_0 = "NO";
    defparam add_1614_17.INJECT1_1 = "NO";
    LUT4 i20020_2_lut (.A(n1025), .B(n1037), .Z(n26708)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i20020_2_lut.init = 16'hdddd;
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (debug_c_c, n30471, GND_net, \register[4] , n13527, 
            n30470, rc_ch4_c, n26947, n1016, n24721, n27035, n30469) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30471;
    input GND_net;
    output [7:0]\register[4] ;
    input n13527;
    input n30470;
    input rc_ch4_c;
    output n26947;
    output n1016;
    input n24721;
    output n27035;
    input n30469;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    wire [15:0]n116;
    
    wire n14954;
    wire [7:0]n43;
    
    wire n4, n4_adj_47, n28543, n28498, n12533, n28467, n28544, 
        n28545, n26527, n28499, n28546, n26475, n24072;
    wire [7:0]n926;
    
    wire n24071, n24070, n24069, n1022, n1010, n26522, n26786, 
        n28398, n26525, n4_adj_48, n28520, n24925, n24719, n26731, 
        n26565, n26315, n54, n19758, n26794, n26067, n24881, n24892, 
        n25, n10, n24028, n24027, n24026, n24025, n24024, n24023, 
        n24022, n24021, n24, n24833, n6, n12141;
    
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_47)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_422 (.A(count[11]), .B(count[10]), .Z(n28543)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_422.init = 16'heeee;
    LUT4 i1_2_lut_rep_377_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n28498)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_377_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_346_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n12533), 
         .D(count[9]), .Z(n28467)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_346_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_423 (.A(count[15]), .B(count[14]), .Z(n28544)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_423.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .D(count[13]), .Z(n12533)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_424 (.A(count[6]), .B(count[7]), .Z(n28545)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_424.init = 16'h8888;
    LUT4 i1_2_lut_rep_378_3_lut (.A(count[6]), .B(count[7]), .C(n26527), 
         .Z(n28499)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_378_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_425 (.A(count[4]), .B(count[5]), .Z(n28546)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_425.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[8]), 
         .D(count[0]), .Z(n26475)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D sub_57_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24072), 
          .S0(n926[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_57_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_9.INIT1 = 16'h0000;
    defparam sub_57_add_2_9.INJECT1_0 = "NO";
    defparam sub_57_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24071), 
          .COUT(n24072), .S0(n926[5]), .S1(n926[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_57_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_7.INJECT1_0 = "NO";
    defparam sub_57_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24070), 
          .COUT(n24071), .S0(n926[3]), .S1(n926[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_57_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_5.INJECT1_0 = "NO";
    defparam sub_57_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24069), 
          .COUT(n24070), .S0(n926[1]), .S1(n926[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_57_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_3.INJECT1_0 = "NO";
    defparam sub_57_add_2_3.INJECT1_1 = "NO";
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n30470), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1022));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1022), .SP(n30470), .CK(debug_c_c), .Q(n1010));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D sub_57_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24069), 
          .S1(n926[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_57_add_2_1.INIT0 = 16'hF000;
    defparam sub_57_add_2_1.INIT1 = 16'h5555;
    defparam sub_57_add_2_1.INJECT1_0 = "NO";
    defparam sub_57_add_2_1.INJECT1_1 = "NO";
    LUT4 count_8__bdd_4_lut (.A(count[8]), .B(n26522), .C(n26786), .D(count[9]), 
         .Z(n28398)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam count_8__bdd_4_lut.init = 16'hf0ee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.A(n26527), .B(n28545), .C(n28546), 
         .D(count[0]), .Z(n26525)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_34.init = 16'h8000;
    LUT4 i1_2_lut (.A(n4_adj_48), .B(n926[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_adj_35 (.A(n4_adj_48), .B(n926[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_35.init = 16'h4444;
    LUT4 i20348_4_lut (.A(n28544), .B(n28520), .C(n24925), .D(n24719), 
         .Z(n26947)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i20348_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n26731), .B(n26565), .C(n28543), .D(n26315), .Z(n24719)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 i3_4_lut (.A(n54), .B(n12533), .C(n4_adj_48), .D(n19758), .Z(n26315)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_36 (.A(n4_adj_48), .B(n926[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_36.init = 16'h4444;
    LUT4 i2_2_lut (.A(n28398), .B(n26794), .Z(n26067)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i2_2_lut.init = 16'h2222;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n24881), .D(n28498), 
         .Z(n24925)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i2_4_lut_adj_37 (.A(n28545), .B(count[5]), .C(count[8]), .D(n4_adj_47), 
         .Z(n24881)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_37.init = 16'ha080;
    LUT4 i5_2_lut_rep_399 (.A(n1010), .B(n1022), .Z(n28520)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_399.init = 16'h4444;
    LUT4 i2_3_lut_4_lut_adj_38 (.A(n1010), .B(n1022), .C(n24925), .D(n28544), 
         .Z(n24892)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i2_3_lut_4_lut_adj_38.init = 16'hfff4;
    LUT4 i20367_4_lut (.A(count[8]), .B(count[7]), .C(n25), .D(count[6]), 
         .Z(n26786)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i20367_4_lut.init = 16'h0001;
    LUT4 i10_3_lut_4_lut (.A(count[8]), .B(n28467), .C(n26525), .D(n26522), 
         .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(160[28:39])
    defparam i10_3_lut_4_lut.init = 16'h0100;
    LUT4 i20039_3_lut_4_lut (.A(count[8]), .B(n28467), .C(n26522), .D(n26525), 
         .Z(n26731)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(160[28:39])
    defparam i20039_3_lut_4_lut.init = 16'hfeee;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    CCU2D add_1610_17 (.A0(count[15]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24028), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_17.INIT0 = 16'hd222;
    defparam add_1610_17.INIT1 = 16'h0000;
    defparam add_1610_17.INJECT1_0 = "NO";
    defparam add_1610_17.INJECT1_1 = "NO";
    CCU2D add_1610_15 (.A0(count[13]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n28520), .C1(GND_net), .D1(GND_net), .CIN(n24027), 
          .COUT(n24028), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_15.INIT0 = 16'hd222;
    defparam add_1610_15.INIT1 = 16'hd222;
    defparam add_1610_15.INJECT1_0 = "NO";
    defparam add_1610_15.INJECT1_1 = "NO";
    CCU2D add_1610_13 (.A0(count[11]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n28520), .C1(GND_net), .D1(GND_net), .CIN(n24026), 
          .COUT(n24027), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_13.INIT0 = 16'hd222;
    defparam add_1610_13.INIT1 = 16'hd222;
    defparam add_1610_13.INJECT1_0 = "NO";
    defparam add_1610_13.INJECT1_1 = "NO";
    CCU2D add_1610_11 (.A0(count[9]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n28520), .C1(GND_net), .D1(GND_net), .CIN(n24025), 
          .COUT(n24026), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_11.INIT0 = 16'hd222;
    defparam add_1610_11.INIT1 = 16'hd222;
    defparam add_1610_11.INJECT1_0 = "NO";
    defparam add_1610_11.INJECT1_1 = "NO";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13527), .PD(n14954), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1610_9 (.A0(count[7]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n28520), .C1(GND_net), .D1(GND_net), .CIN(n24024), 
          .COUT(n24025), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_9.INIT0 = 16'hd222;
    defparam add_1610_9.INIT1 = 16'hd222;
    defparam add_1610_9.INJECT1_0 = "NO";
    defparam add_1610_9.INJECT1_1 = "NO";
    CCU2D add_1610_7 (.A0(count[5]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n28520), .C1(GND_net), .D1(GND_net), .CIN(n24023), 
          .COUT(n24024), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_7.INIT0 = 16'hd222;
    defparam add_1610_7.INIT1 = 16'hd222;
    defparam add_1610_7.INJECT1_0 = "NO";
    defparam add_1610_7.INJECT1_1 = "NO";
    CCU2D add_1610_5 (.A0(count[3]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n28520), .C1(GND_net), .D1(GND_net), .CIN(n24022), 
          .COUT(n24023), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_5.INIT0 = 16'hd222;
    defparam add_1610_5.INIT1 = 16'hd222;
    defparam add_1610_5.INJECT1_0 = "NO";
    defparam add_1610_5.INJECT1_1 = "NO";
    CCU2D add_1610_3 (.A0(count[1]), .B0(n28520), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n28520), .C1(GND_net), .D1(GND_net), .CIN(n24021), 
          .COUT(n24022), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_3.INIT0 = 16'hd222;
    defparam add_1610_3.INIT1 = 16'hd222;
    defparam add_1610_3.INJECT1_0 = "NO";
    defparam add_1610_3.INJECT1_1 = "NO";
    FD1P3AX valid_48 (.D(n26067), .SP(n24721), .CK(debug_c_c), .Q(n1016));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D add_1610_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n24892), .B1(n1022), .C1(count[0]), .D1(n1010), .COUT(n24021), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1610_1.INIT0 = 16'hF000;
    defparam add_1610_1.INIT1 = 16'ha565;
    defparam add_1610_1.INJECT1_0 = "NO";
    defparam add_1610_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_39 (.A(n4_adj_48), .B(n926[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_39.init = 16'h4444;
    LUT4 i20436_4_lut (.A(n54), .B(n26565), .C(n4_adj_48), .D(n10), 
         .Z(n27035)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i20436_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_40 (.A(n30469), .B(n26794), .C(n24), .D(n26565), 
         .Z(n14954)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_40.init = 16'h0020;
    LUT4 i31_4_lut (.A(n28499), .B(n24833), .C(count[9]), .D(n26475), 
         .Z(n24)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_4_lut.init = 16'h3a30;
    LUT4 i1_2_lut_adj_41 (.A(n4_adj_48), .B(n926[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_41.init = 16'h4444;
    LUT4 i2_4_lut_adj_42 (.A(n28499), .B(n28467), .C(n28546), .D(count[8]), 
         .Z(n4_adj_48)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_42.init = 16'hecff;
    LUT4 i3_4_lut_adj_43 (.A(n25), .B(count[6]), .C(count[8]), .D(count[7]), 
         .Z(n24833)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_43.init = 16'hfffe;
    LUT4 i1_4_lut_adj_44 (.A(count[0]), .B(n28546), .C(n6), .D(count[3]), 
         .Z(n25)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_44.init = 16'hccc8;
    LUT4 i2_2_lut_adj_45 (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_45.init = 16'heeee;
    LUT4 i2_3_lut (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n26527)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i20098_4_lut (.A(count[12]), .B(n28544), .C(count[13]), .D(n28543), 
         .Z(n26794)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20098_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_46 (.A(n1022), .B(n1010), .Z(n26565)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_46.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_47 (.A(n28545), .B(count[5]), .C(count[4]), .D(n4), 
         .Z(n26522)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_47.init = 16'h8880;
    LUT4 i21_4_lut (.A(n12141), .B(n12533), .C(n19758), .D(n28543), 
         .Z(n54)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h0002;
    LUT4 i1_4_lut_adj_48 (.A(n26475), .B(n28467), .C(n28545), .D(n26527), 
         .Z(n12141)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_48.init = 16'heccc;
    LUT4 i13777_2_lut (.A(n24833), .B(count[9]), .Z(n19758)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13777_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_49 (.A(n4_adj_48), .B(n926[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_49.init = 16'h4444;
    LUT4 i1_2_lut_adj_50 (.A(n4_adj_48), .B(n926[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_50.init = 16'h4444;
    LUT4 i1_2_lut_adj_51 (.A(n4_adj_48), .B(n926[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_51.init = 16'h4444;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (debug_c_c, n30471, GND_net, \register[3] , n13534, 
            n30470, rc_ch3_c, n27027, n30469, n26939, n1001, n24755) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30471;
    input GND_net;
    output [7:0]\register[3] ;
    input n13534;
    input n30470;
    input rc_ch3_c;
    output n27027;
    input n30469;
    output n26939;
    output n1001;
    input n24755;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    wire [15:0]n116;
    
    wire n14957;
    wire [7:0]n43;
    
    wire n995, n1007, n28533, n24926, n28572, n26605, n28512, 
        n24076;
    wire [7:0]n917;
    
    wire n24075, n24074, n24073, n28478, n26539, n24610, n10, 
        n26719, n28513, n28479, n12441, n28424, n26760, n26537, 
        n28423, n28450, n26606, n28552, n28569, n103, n5, n28571, 
        n4, n28573, n4_adj_45, n26778, n28570, n152, n154, n26589, 
        n11, n24754, n24036, n24035, n24034, n24033, n4_adj_46, 
        n24032, n24031, n24030, n24029, n6;
    
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    LUT4 i5_2_lut_rep_412 (.A(n995), .B(n1007), .Z(n28533)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_412.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n995), .B(n1007), .C(n24926), .D(n28572), 
         .Z(n26605)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_rep_391_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n28512)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_391_3_lut.init = 16'h8080;
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D sub_56_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24076), 
          .S0(n917[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_56_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_9.INIT1 = 16'h0000;
    defparam sub_56_add_2_9.INJECT1_0 = "NO";
    defparam sub_56_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24075), 
          .COUT(n24076), .S0(n917[5]), .S1(n917[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_56_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_7.INJECT1_0 = "NO";
    defparam sub_56_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24074), 
          .COUT(n24075), .S0(n917[3]), .S1(n917[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_56_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_5.INJECT1_0 = "NO";
    defparam sub_56_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24073), 
          .COUT(n24074), .S0(n917[1]), .S1(n917[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_56_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_3.INJECT1_0 = "NO";
    defparam sub_56_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24073), 
          .S1(n917[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_56_add_2_1.INIT0 = 16'hF000;
    defparam sub_56_add_2_1.INIT1 = 16'h5555;
    defparam sub_56_add_2_1.INJECT1_0 = "NO";
    defparam sub_56_add_2_1.INJECT1_1 = "NO";
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n28478), .C(n26539), 
         .D(n24610), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i20030_3_lut_4_lut (.A(count[8]), .B(n28478), .C(n24610), .D(n26539), 
         .Z(n26719)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i20030_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_28 (.A(count[7]), .B(count[6]), .C(count[0]), 
         .D(n28513), .Z(n26539)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut_adj_28.init = 16'h8000;
    LUT4 i13675_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13675_2_lut_4_lut.init = 16'h0400;
    LUT4 i13674_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13674_2_lut_4_lut.init = 16'h0400;
    LUT4 i13673_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13673_2_lut_4_lut.init = 16'h0400;
    LUT4 i13672_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13672_2_lut_4_lut.init = 16'h0400;
    LUT4 i13671_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13671_2_lut_4_lut.init = 16'h0400;
    LUT4 i13670_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13670_2_lut_4_lut.init = 16'h0400;
    LUT4 i13669_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13669_2_lut_4_lut.init = 16'h0400;
    LUT4 i13455_2_lut_4_lut (.A(n28478), .B(count[8]), .C(n28479), .D(n917[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13455_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_357 (.A(count[9]), .B(n12441), .Z(n28478)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_357.init = 16'heeee;
    LUT4 i1_2_lut_rep_303_3_lut_4_lut (.A(count[9]), .B(n12441), .C(n24610), 
         .D(count[8]), .Z(n28424)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_303_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21_3_lut_rep_302_4_lut (.A(count[9]), .B(n12441), .C(n26760), 
         .D(n26537), .Z(n28423)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i21_3_lut_rep_302_4_lut.init = 16'h0f0e;
    LUT4 i1_3_lut_rep_329_4_lut (.A(count[9]), .B(n12441), .C(n28479), 
         .D(count[8]), .Z(n28450)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_3_lut_rep_329_4_lut.init = 16'hfeff;
    LUT4 i20382_3_lut_3_lut_4_lut (.A(n28572), .B(n24926), .C(n28424), 
         .D(n26760), .Z(n26606)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i20382_3_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3AX prev_in_46 (.D(n1007), .SP(n30470), .CK(debug_c_c), .Q(n995));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n30470), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1007));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_431 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n28552)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_431.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[8]), .D(n28569), 
         .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_451 (.A(count[15]), .B(count[14]), .Z(n28572)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_451.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_29 (.A(n26537), .B(n26760), .C(n28478), .D(n28450), 
         .Z(n5)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut_adj_29.init = 16'hcd00;
    LUT4 i1_2_lut_rep_450 (.A(count[7]), .B(count[6]), .Z(n28571)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_450.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_452 (.A(count[11]), .B(count[10]), .Z(n28573)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_452.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4_adj_45)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i20084_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n26778)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20084_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_449 (.A(count[2]), .B(count[1]), .Z(n28570)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_449.init = 16'h8888;
    LUT4 i2_3_lut_rep_392_4_lut (.A(count[4]), .B(count[5]), .C(n28570), 
         .D(count[3]), .Z(n28513)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_rep_392_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_448 (.A(count[4]), .B(count[5]), .Z(n28569)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_448.init = 16'h8888;
    PFUMX i12645 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    LUT4 i20428_4_lut (.A(n28423), .B(n26589), .C(n28450), .D(n10), 
         .Z(n27027)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i20428_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n30469), .B(n28572), .C(n11), .D(n26778), .Z(n14957)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i4_4_lut (.A(n26537), .B(n26589), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i1_3_lut_4_lut_adj_30 (.A(count[8]), .B(n28571), .C(count[0]), 
         .D(n28513), .Z(n26537)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_4_lut_adj_30.init = 16'h8000;
    LUT4 i1_2_lut_rep_358_4_lut (.A(count[3]), .B(n28570), .C(n28569), 
         .D(n28571), .Z(n28479)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_358_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(n1007), .B(n995), .Z(n26589)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i20340_4_lut (.A(n28572), .B(n28533), .C(n24926), .D(n24754), 
         .Z(n26939)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i20340_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5), .B(n26589), .C(n26719), .D(n26760), .Z(n24754)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i2_4_lut_adj_31 (.A(n28571), .B(count[5]), .C(count[3]), .D(n4_adj_45), 
         .Z(n24610)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_31.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n28572), .D(n28573), 
         .Z(n12441)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i20066_3_lut (.A(n12441), .B(count[9]), .C(n154), .Z(n26760)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i20066_3_lut.init = 16'heaea;
    CCU2D add_1606_17 (.A0(count[15]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24036), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_17.INIT0 = 16'hd222;
    defparam add_1606_17.INIT1 = 16'h0000;
    defparam add_1606_17.INJECT1_0 = "NO";
    defparam add_1606_17.INJECT1_1 = "NO";
    CCU2D add_1606_15 (.A0(count[13]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n28533), .C1(GND_net), .D1(GND_net), .CIN(n24035), 
          .COUT(n24036), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_15.INIT0 = 16'hd222;
    defparam add_1606_15.INIT1 = 16'hd222;
    defparam add_1606_15.INJECT1_0 = "NO";
    defparam add_1606_15.INJECT1_1 = "NO";
    CCU2D add_1606_13 (.A0(count[11]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n28533), .C1(GND_net), .D1(GND_net), .CIN(n24034), 
          .COUT(n24035), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_13.INIT0 = 16'hd222;
    defparam add_1606_13.INIT1 = 16'hd222;
    defparam add_1606_13.INJECT1_0 = "NO";
    defparam add_1606_13.INJECT1_1 = "NO";
    CCU2D add_1606_11 (.A0(count[9]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n28533), .C1(GND_net), .D1(GND_net), .CIN(n24033), 
          .COUT(n24034), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_11.INIT0 = 16'hd222;
    defparam add_1606_11.INIT1 = 16'hd222;
    defparam add_1606_11.INJECT1_0 = "NO";
    defparam add_1606_11.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_32 (.A(count[13]), .B(count[12]), .C(n28573), .D(n4_adj_46), 
         .Z(n24926)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_32.init = 16'h8880;
    CCU2D add_1606_9 (.A0(count[7]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n28533), .C1(GND_net), .D1(GND_net), .CIN(n24032), 
          .COUT(n24033), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_9.INIT0 = 16'hd222;
    defparam add_1606_9.INIT1 = 16'hd222;
    defparam add_1606_9.INJECT1_0 = "NO";
    defparam add_1606_9.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13534), .PD(n14957), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1606_7 (.A0(count[5]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n28533), .C1(GND_net), .D1(GND_net), .CIN(n24031), 
          .COUT(n24032), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_7.INIT0 = 16'hd222;
    defparam add_1606_7.INIT1 = 16'hd222;
    defparam add_1606_7.INJECT1_0 = "NO";
    defparam add_1606_7.INJECT1_1 = "NO";
    CCU2D add_1606_5 (.A0(count[3]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n28533), .C1(GND_net), .D1(GND_net), .CIN(n24030), 
          .COUT(n24031), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_5.INIT0 = 16'hd222;
    defparam add_1606_5.INIT1 = 16'hd222;
    defparam add_1606_5.INJECT1_0 = "NO";
    defparam add_1606_5.INJECT1_1 = "NO";
    CCU2D add_1606_3 (.A0(count[1]), .B0(n28533), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n28533), .C1(GND_net), .D1(GND_net), .CIN(n24029), 
          .COUT(n24030), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_3.INIT0 = 16'hd222;
    defparam add_1606_3.INIT1 = 16'hd222;
    defparam add_1606_3.INJECT1_0 = "NO";
    defparam add_1606_3.INJECT1_1 = "NO";
    LUT4 i23_4_lut (.A(n28552), .B(count[2]), .C(n28569), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    CCU2D add_1606_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n26605), .B1(n1007), .C1(count[0]), .D1(n995), .COUT(n24029), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1606_1.INIT0 = 16'hF000;
    defparam add_1606_1.INIT1 = 16'ha565;
    defparam add_1606_1.INJECT1_0 = "NO";
    defparam add_1606_1.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_33 (.A(count[9]), .B(count[4]), .C(n28512), .D(n4), 
         .Z(n4_adj_46)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_33.init = 16'hfaea;
    FD1P3IX valid_48 (.D(n26606), .SP(n24755), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1001));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (GND_net, debug_c_c, n30470, rc_ch2_c, n26945, 
            \register[2] , n13535, n986, n24741, n27025, n30469, 
            n28403, n30471) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n30470;
    input rc_ch2_c;
    output n26945;
    output [7:0]\register[2] ;
    input n13535;
    output n986;
    input n24741;
    output n27025;
    input n30469;
    input n28403;
    input n30471;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24078;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    wire [7:0]n908;
    
    wire n24079, n24077, n28463, n28436, n24582, n10, n26723, 
        n28462;
    wire [7:0]n43;
    
    wire n28538, n28495, n28539, n6, n4, n54, n5, n4_adj_40, 
        n28540, n26776, n28541, n24927, n28418, n5_adj_41, n26614, 
        n992, n28550, n28551, n103, n28491, n5_adj_42, n28434, 
        n26752, n26615, n152, n154, n24044;
    wire [15:0]n116;
    
    wire n24043, n24042, n24041, n24740, n26712, n24040, n24039, 
        n24038, n24037, n980, n26534, n4_adj_43, n14959, n6_adj_44, 
        n12412, n28435, n11, n24080;
    
    CCU2D sub_55_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24078), 
          .COUT(n24079), .S0(n908[3]), .S1(n908[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_55_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_55_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_55_add_2_5.INJECT1_0 = "NO";
    defparam sub_55_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_55_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24077), 
          .COUT(n24078), .S0(n908[1]), .S1(n908[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_55_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_55_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_55_add_2_3.INJECT1_0 = "NO";
    defparam sub_55_add_2_3.INJECT1_1 = "NO";
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n28463), .C(n28436), 
         .D(n24582), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    CCU2D sub_55_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24077), 
          .S1(n908[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_55_add_2_1.INIT0 = 16'hF000;
    defparam sub_55_add_2_1.INIT1 = 16'h5555;
    defparam sub_55_add_2_1.INJECT1_0 = "NO";
    defparam sub_55_add_2_1.INJECT1_1 = "NO";
    LUT4 i20032_3_lut_4_lut (.A(count[8]), .B(n28463), .C(n24582), .D(n28436), 
         .Z(n26723)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i20032_3_lut_4_lut.init = 16'hfeee;
    LUT4 i13442_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13442_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_417 (.A(count[7]), .B(count[6]), .Z(n28538)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_417.init = 16'h8888;
    LUT4 i1_2_lut_rep_374_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n28495)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_374_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n28539), 
         .D(count[8]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_418 (.A(count[2]), .B(count[1]), .Z(n28539)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_418.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n54), 
         .Z(n5)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h00fb;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4_adj_40)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i13666_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13666_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_419 (.A(count[10]), .B(count[11]), .Z(n28540)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_419.init = 16'heeee;
    LUT4 i20082_3_lut_4_lut (.A(count[10]), .B(count[11]), .C(count[13]), 
         .D(count[12]), .Z(n26776)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20082_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_420 (.A(count[15]), .B(count[14]), .Z(n28541)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_420.init = 16'heeee;
    LUT4 i1_2_lut_rep_297_3_lut (.A(count[15]), .B(count[14]), .C(n24927), 
         .Z(n28418)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_297_3_lut.init = 16'hfefe;
    LUT4 i13665_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13665_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5_adj_41), 
         .D(n24927), .Z(n26614)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i13664_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13664_2_lut_4_lut.init = 16'h0400;
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n30470), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n992));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_429 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n28550)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_429.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_22 (.A(count[7]), .B(count[6]), .C(count[8]), 
         .D(n28551), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_22.init = 16'hfffe;
    LUT4 i1_2_lut_rep_430 (.A(count[4]), .B(count[5]), .Z(n28551)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_430.init = 16'h8888;
    LUT4 i1_2_lut_rep_370_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n28491)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_370_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n5_adj_42)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut_adj_23.init = 16'h8000;
    LUT4 i13663_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13663_2_lut_4_lut.init = 16'h0400;
    LUT4 i13662_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13662_2_lut_4_lut.init = 16'h0400;
    LUT4 i20380_3_lut_3_lut_4_lut (.A(n24582), .B(n28434), .C(n26752), 
         .D(n28418), .Z(n26615)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i20380_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i3_3_lut_rep_341_4_lut (.A(count[3]), .B(n28551), .C(n28538), 
         .D(n28539), .Z(n28462)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_3_lut_rep_341_4_lut.init = 16'h8000;
    LUT4 i13661_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13661_2_lut_4_lut.init = 16'h0400;
    PFUMX i12739 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    CCU2D add_1602_17 (.A0(count[15]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24044), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_17.INIT0 = 16'hd222;
    defparam add_1602_17.INIT1 = 16'h0000;
    defparam add_1602_17.INJECT1_0 = "NO";
    defparam add_1602_17.INJECT1_1 = "NO";
    CCU2D add_1602_15 (.A0(count[13]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5_adj_41), .C1(GND_net), .D1(GND_net), 
          .CIN(n24043), .COUT(n24044), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_15.INIT0 = 16'hd222;
    defparam add_1602_15.INIT1 = 16'hd222;
    defparam add_1602_15.INJECT1_0 = "NO";
    defparam add_1602_15.INJECT1_1 = "NO";
    CCU2D add_1602_13 (.A0(count[11]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5_adj_41), .C1(GND_net), .D1(GND_net), 
          .CIN(n24042), .COUT(n24043), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_13.INIT0 = 16'hd222;
    defparam add_1602_13.INIT1 = 16'hd222;
    defparam add_1602_13.INJECT1_0 = "NO";
    defparam add_1602_13.INJECT1_1 = "NO";
    CCU2D add_1602_11 (.A0(count[9]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5_adj_41), .C1(GND_net), .D1(GND_net), 
          .CIN(n24041), .COUT(n24042), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_11.INIT0 = 16'hd222;
    defparam add_1602_11.INIT1 = 16'hd222;
    defparam add_1602_11.INJECT1_0 = "NO";
    defparam add_1602_11.INJECT1_1 = "NO";
    LUT4 i20346_4_lut (.A(n28541), .B(n5_adj_41), .C(n24927), .D(n24740), 
         .Z(n26945)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i20346_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5), .B(n26712), .C(n26723), .D(n26752), .Z(n24740)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    CCU2D add_1602_9 (.A0(count[7]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5_adj_41), .C1(GND_net), .D1(GND_net), 
          .CIN(n24040), .COUT(n24041), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_9.INIT0 = 16'hd222;
    defparam add_1602_9.INIT1 = 16'hd222;
    defparam add_1602_9.INJECT1_0 = "NO";
    defparam add_1602_9.INJECT1_1 = "NO";
    CCU2D add_1602_7 (.A0(count[5]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5_adj_41), .C1(GND_net), .D1(GND_net), 
          .CIN(n24039), .COUT(n24040), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_7.INIT0 = 16'hd222;
    defparam add_1602_7.INIT1 = 16'hd222;
    defparam add_1602_7.INJECT1_0 = "NO";
    defparam add_1602_7.INJECT1_1 = "NO";
    CCU2D add_1602_5 (.A0(count[3]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5_adj_41), .C1(GND_net), .D1(GND_net), 
          .CIN(n24038), .COUT(n24039), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_5.INIT0 = 16'hd222;
    defparam add_1602_5.INIT1 = 16'hd222;
    defparam add_1602_5.INJECT1_0 = "NO";
    defparam add_1602_5.INJECT1_1 = "NO";
    CCU2D add_1602_3 (.A0(count[1]), .B0(n5_adj_41), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5_adj_41), .C1(GND_net), .D1(GND_net), 
          .CIN(n24037), .COUT(n24038), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_3.INIT0 = 16'hd222;
    defparam add_1602_3.INIT1 = 16'hd222;
    defparam add_1602_3.INJECT1_0 = "NO";
    defparam add_1602_3.INJECT1_1 = "NO";
    CCU2D add_1602_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n26614), .B1(n992), .C1(count[0]), .D1(n980), .COUT(n24037), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1602_1.INIT0 = 16'hF000;
    defparam add_1602_1.INIT1 = 16'ha565;
    defparam add_1602_1.INJECT1_0 = "NO";
    defparam add_1602_1.INJECT1_1 = "NO";
    LUT4 i13660_2_lut_4_lut (.A(n28463), .B(count[8]), .C(n28462), .D(n908[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i13660_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_adj_24 (.A(count[0]), .B(n28462), .C(count[8]), 
         .Z(n26534)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_24.init = 16'h8080;
    FD1P3AX prev_in_46 (.D(n992), .SP(n30470), .CK(debug_c_c), .Q(n980));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n28540), .D(n4_adj_43), 
         .Z(n24927)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i23_4_lut (.A(n28550), .B(count[2]), .C(n28551), .D(n6_adj_44), 
         .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6_adj_44)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_25 (.A(count[9]), .B(count[4]), .C(n28495), .D(n4_adj_40), 
         .Z(n4_adj_43)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_25.init = 16'hfaea;
    FD1P3IX valid_48 (.D(n26615), .SP(n24741), .CD(GND_net), .CK(debug_c_c), 
            .Q(n986));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_315_4_lut (.A(n28539), .B(n28538), .C(n28491), .D(count[0]), 
         .Z(n28436)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_315_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_342 (.A(count[9]), .B(n12412), .Z(n28463)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_342.init = 16'heeee;
    LUT4 i1_2_lut_rep_313_3_lut (.A(count[9]), .B(n12412), .C(count[8]), 
         .Z(n28434)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_313_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_rep_314_4_lut (.A(count[9]), .B(n12412), .C(n28462), 
         .D(count[8]), .Z(n28435)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_3_lut_rep_314_4_lut.init = 16'hfeff;
    LUT4 i5_2_lut (.A(n980), .B(n992), .Z(n5_adj_41)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i20426_4_lut (.A(n54), .B(n26712), .C(n28435), .D(n10), .Z(n27025)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i20426_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_26 (.A(n30469), .B(n28541), .C(n11), .D(n26776), 
         .Z(n14959)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_26.init = 16'h0020;
    LUT4 i4_4_lut (.A(n26534), .B(n26712), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n28541), .D(n28540), 
         .Z(n12412)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i20024_2_lut (.A(n980), .B(n992), .Z(n26712)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i20024_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_adj_27 (.A(n28538), .B(count[5]), .C(count[3]), .D(n4), 
         .Z(n24582)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_27.init = 16'h8880;
    LUT4 i21_4_lut (.A(n5_adj_42), .B(n26752), .C(n28463), .D(n6), .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i20058_3_lut (.A(n12412), .B(count[9]), .C(n154), .Z(n26752)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i20058_3_lut.init = 16'heaea;
    CCU2D sub_55_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24080), 
          .S0(n908[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_55_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_55_add_2_9.INIT1 = 16'h0000;
    defparam sub_55_add_2_9.INJECT1_0 = "NO";
    defparam sub_55_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_55_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24079), 
          .COUT(n24080), .S0(n908[5]), .S1(n908[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_55_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_55_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_55_add_2_7.INJECT1_0 = "NO";
    defparam sub_55_add_2_7.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n28403), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n28403), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n28403), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n28403), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n28403), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n28403), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n28403), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n28403), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30471), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30471), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13535), .PD(n14959), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (debug_c_c, n30470, n26907, rc_ch1_c, GND_net, 
            \register[1] , n13536, n971, n24716, n27023, n30469) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30470;
    output n26907;
    input rc_ch1_c;
    input GND_net;
    output [7:0]\register[1] ;
    input n13536;
    output n971;
    input n24716;
    output n27023;
    input n30469;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n4, n4_adj_39, n28529, n28492, n12539, n28465, n28530, 
        n5, n24928, n26597, n28429, n28531, n26466, n28493, n28532, 
        n28494, n965, n977, n24713, n26733, n26607, n26313, n54, 
        n26290, n28464, n24878, n24529, n28437, n24899, n26596, 
        n26458;
    wire [7:0]n899;
    wire [7:0]n43;
    
    wire n10;
    wire [15:0]n116;
    
    wire n14962, n26343, n24, n26531, n24826, n24794, n6, n24448, 
        n24447, n24446, n24445, n24444, n24443, n24442, n24441, 
        n24084, n24083, n24082, n24081;
    
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_39)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_408 (.A(count[11]), .B(count[10]), .Z(n28529)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_408.init = 16'heeee;
    LUT4 i1_2_lut_rep_371_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n28492)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_371_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n12539), 
         .D(count[9]), .Z(n28465)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_409 (.A(count[15]), .B(count[14]), .Z(n28530)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_409.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n12539)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n24928), 
         .Z(n26597)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_308_3_lut (.A(count[15]), .B(count[14]), .C(n24928), 
         .Z(n28429)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_308_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_410 (.A(count[6]), .B(count[7]), .Z(n28531)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_410.init = 16'h8888;
    LUT4 i1_2_lut_rep_372_3_lut (.A(count[6]), .B(count[7]), .C(n26466), 
         .Z(n28493)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_372_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_411 (.A(count[4]), .B(count[5]), .Z(n28532)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_411.init = 16'h8888;
    LUT4 i1_2_lut_rep_373_3_lut (.A(count[4]), .B(count[5]), .C(count[0]), 
         .Z(n28494)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_373_3_lut.init = 16'h8080;
    FD1P3AX prev_in_46 (.D(n977), .SP(n30470), .CK(debug_c_c), .Q(n965));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i20308_4_lut (.A(n28530), .B(n5), .C(n24928), .D(n24713), .Z(n26907)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i20308_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n26733), .B(n26607), .C(n28529), .D(n26313), .Z(n24713)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 i3_4_lut (.A(n54), .B(n12539), .C(n26290), .D(n28464), .Z(n26313)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i5_2_lut (.A(n965), .B(n977), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n24878), .D(n28492), 
         .Z(n24928)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i2_4_lut_adj_5 (.A(n28531), .B(count[5]), .C(count[8]), .D(n4_adj_39), 
         .Z(n24878)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_5.init = 16'ha080;
    LUT4 i20312_3_lut_3_lut_4_lut (.A(n24529), .B(n28437), .C(n24899), 
         .D(n28429), .Z(n26596)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i20312_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_2_lut_rep_316_3_lut_4_lut (.A(count[9]), .B(n28529), .C(count[8]), 
         .D(n12539), .Z(n28437)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_316_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_6 (.A(count[0]), .B(n28532), .C(n28531), 
         .D(n26466), .Z(n26458)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_6.init = 16'h8000;
    LUT4 i1_2_lut (.A(n26290), .B(n899[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_adj_7 (.A(n26290), .B(n899[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_7.init = 16'h4444;
    LUT4 i1_2_lut_adj_8 (.A(n26290), .B(n899[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_8.init = 16'h4444;
    LUT4 i1_2_lut_adj_9 (.A(n26290), .B(n899[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_9.init = 16'h4444;
    LUT4 i1_2_lut_adj_10 (.A(n26290), .B(n899[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_10.init = 16'h4444;
    LUT4 i1_2_lut_adj_11 (.A(n26290), .B(n899[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_11.init = 16'h4444;
    LUT4 i1_2_lut_adj_12 (.A(n26290), .B(n899[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_12.init = 16'h4444;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n28465), .C(n26458), 
         .D(n24529), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i20040_3_lut_4_lut (.A(count[8]), .B(n28465), .C(n24529), .D(n26458), 
         .Z(n26733)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i20040_3_lut_4_lut.init = 16'hfeee;
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n30470), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n977));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3AX valid_48 (.D(n26596), .SP(n24716), .CK(debug_c_c), .Q(n971));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    LUT4 i20424_4_lut (.A(n54), .B(n26607), .C(n26290), .D(n10), .Z(n27023)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i20424_4_lut.init = 16'h3323;
    LUT4 i3_4_lut_adj_13 (.A(n28530), .B(n26343), .C(n28529), .D(n30469), 
         .Z(n14962)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_13.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[13]), .B(n24), .C(count[12]), .D(n26607), 
         .Z(n26343)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i31_3_lut (.A(n26531), .B(n24826), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30470), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_14 (.A(n26290), .B(n899[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_14.init = 16'h4444;
    LUT4 i1_4_lut_adj_15 (.A(n28465), .B(count[8]), .C(n28493), .D(n28532), 
         .Z(n26290)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_15.init = 16'hfbbb;
    LUT4 i1_4_lut_adj_16 (.A(n26466), .B(n28531), .C(count[8]), .D(n28494), 
         .Z(n26531)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_16.init = 16'h8000;
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30470), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_17 (.A(n24794), .B(n6), .C(count[8]), .D(n28532), 
         .Z(n24826)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_17.init = 16'hfefc;
    LUT4 i3_4_lut_adj_18 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n24794)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_18.init = 16'hfffe;
    LUT4 i13775_2_lut_rep_343 (.A(n24826), .B(count[9]), .Z(n28464)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13775_2_lut_rep_343.init = 16'h8888;
    LUT4 i2_3_lut_4_lut_adj_19 (.A(n24826), .B(count[9]), .C(n28529), 
         .D(n12539), .Z(n24899)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i2_3_lut_4_lut_adj_19.init = 16'hfff8;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n26466)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_adj_20 (.A(n977), .B(n965), .Z(n26607)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_20.init = 16'hbbbb;
    CCU2D add_1598_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24448), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_17.INIT0 = 16'hd222;
    defparam add_1598_17.INIT1 = 16'h0000;
    defparam add_1598_17.INJECT1_0 = "NO";
    defparam add_1598_17.INJECT1_1 = "NO";
    CCU2D add_1598_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n24447), 
          .COUT(n24448), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_15.INIT0 = 16'hd222;
    defparam add_1598_15.INIT1 = 16'hd222;
    defparam add_1598_15.INJECT1_0 = "NO";
    defparam add_1598_15.INJECT1_1 = "NO";
    CCU2D add_1598_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n24446), 
          .COUT(n24447), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_13.INIT0 = 16'hd222;
    defparam add_1598_13.INIT1 = 16'hd222;
    defparam add_1598_13.INJECT1_0 = "NO";
    defparam add_1598_13.INJECT1_1 = "NO";
    CCU2D add_1598_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n24445), 
          .COUT(n24446), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_11.INIT0 = 16'hd222;
    defparam add_1598_11.INIT1 = 16'hd222;
    defparam add_1598_11.INJECT1_0 = "NO";
    defparam add_1598_11.INJECT1_1 = "NO";
    CCU2D add_1598_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n24444), 
          .COUT(n24445), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_9.INIT0 = 16'hd222;
    defparam add_1598_9.INIT1 = 16'hd222;
    defparam add_1598_9.INJECT1_0 = "NO";
    defparam add_1598_9.INJECT1_1 = "NO";
    LUT4 i21_3_lut_4_lut (.A(n12539), .B(n28492), .C(n24899), .D(n26531), 
         .Z(n54)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i21_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i2_4_lut_adj_21 (.A(n28531), .B(count[4]), .C(count[5]), .D(n4), 
         .Z(n24529)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_21.init = 16'ha080;
    CCU2D add_1598_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n24443), 
          .COUT(n24444), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_7.INIT0 = 16'hd222;
    defparam add_1598_7.INIT1 = 16'hd222;
    defparam add_1598_7.INJECT1_0 = "NO";
    defparam add_1598_7.INJECT1_1 = "NO";
    CCU2D add_1598_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n24442), 
          .COUT(n24443), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_5.INIT0 = 16'hd222;
    defparam add_1598_5.INIT1 = 16'hd222;
    defparam add_1598_5.INJECT1_0 = "NO";
    defparam add_1598_5.INJECT1_1 = "NO";
    CCU2D add_1598_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n24441), 
          .COUT(n24442), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_3.INIT0 = 16'hd222;
    defparam add_1598_3.INIT1 = 16'hd222;
    defparam add_1598_3.INJECT1_0 = "NO";
    defparam add_1598_3.INJECT1_1 = "NO";
    CCU2D add_1598_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n26597), .B1(n977), .C1(count[0]), .D1(n965), .COUT(n24441), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1598_1.INIT0 = 16'hF000;
    defparam add_1598_1.INIT1 = 16'ha565;
    defparam add_1598_1.INJECT1_0 = "NO";
    defparam add_1598_1.INJECT1_1 = "NO";
    CCU2D sub_54_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24084), 
          .S0(n899[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_54_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_54_add_2_9.INIT1 = 16'h0000;
    defparam sub_54_add_2_9.INJECT1_0 = "NO";
    defparam sub_54_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_54_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24083), 
          .COUT(n24084), .S0(n899[5]), .S1(n899[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_54_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_54_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_54_add_2_7.INJECT1_0 = "NO";
    defparam sub_54_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_54_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24082), 
          .COUT(n24083), .S0(n899[3]), .S1(n899[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_54_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_54_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_54_add_2_5.INJECT1_0 = "NO";
    defparam sub_54_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_54_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24081), 
          .COUT(n24082), .S0(n899[1]), .S1(n899[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_54_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_54_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_54_add_2_3.INJECT1_0 = "NO";
    defparam sub_54_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_54_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24081), 
          .S1(n899[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_54_add_2_1.INIT0 = 16'hF000;
    defparam sub_54_add_2_1.INIT1 = 16'h5555;
    defparam sub_54_add_2_1.INJECT1_0 = "NO";
    defparam sub_54_add_2_1.INJECT1_1 = "NO";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13536), .PD(n14962), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (\register_addr[1] , n24822, 
            debug_c_c, VCC_net, GND_net, Stepper_Y_nFault_c, n28477, 
            \read_size[0] , n2622, n26514, Stepper_Y_M0_c_0, n12650, 
            n579, prev_step_clk, step_clk, limit_latched, prev_limit_latched, 
            n13363, prev_select, n28452, read_value, \register_addr[0] , 
            Stepper_Y_M1_c_1, databus, n3539, n32, limit_c_1, Stepper_Y_Dir_c, 
            Stepper_Y_En_c, n8273, n611, \control_reg[7] , n12649, 
            n11054, Stepper_Y_M2_c_2, \read_size[2] , n26540, Stepper_Y_Step_c, 
            n22, n28411, n7685, n28400, n14873, n7244, n7278) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[1] ;
    output n24822;
    input debug_c_c;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    input n28477;
    output \read_size[0] ;
    input n2622;
    input n26514;
    output Stepper_Y_M0_c_0;
    input n12650;
    input n579;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    input n13363;
    output prev_select;
    input n28452;
    output [31:0]read_value;
    input \register_addr[0] ;
    output Stepper_Y_M1_c_1;
    input [31:0]databus;
    input n3539;
    input n32;
    input limit_c_1;
    output Stepper_Y_Dir_c;
    output Stepper_Y_En_c;
    input n8273;
    input n611;
    output \control_reg[7] ;
    input n12649;
    input n11054;
    output Stepper_Y_M2_c_2;
    output \read_size[2] ;
    input n26540;
    output Stepper_Y_Step_c;
    input n22;
    input n28411;
    input n7685;
    input n28400;
    input n14873;
    output n7244;
    output n7278;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n26805, n26806, n26807, n49, n62, n58, n50;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n41, n60, n54, n42, n52, n38, n56, n46, n26823, n26824, 
        n26825, fault_latched;
    wire [31:0]n3540;
    
    wire n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [7:0]n7684;
    wire [31:0]n5671;
    wire [31:0]n100;
    
    wire n26867;
    wire [31:0]n224;
    
    wire n24196, n24195, n24194, n24193, n24192, n24191, n24190, 
        n24189, n24188, n24187, n24186, n24185, n24184, n24183, 
        n24182, n24181, n26865, n26866, int_step;
    
    PFUMX i20111 (.BLUT(n26805), .ALUT(n26806), .C0(\register_addr[1] ), 
          .Z(n26807));
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n24822)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(steps_reg[9]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(steps_reg[3]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    PFUMX i20129 (.BLUT(n26823), .ALUT(n26824), .C0(\register_addr[1] ), 
          .Z(n26825));
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[6]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3540[0]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n26514), .SP(n2622), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12650), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13363), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n28452), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n26807), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i13255_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7684[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13255_2_lut.init = 16'h2222;
    LUT4 mux_1755_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5671[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1755_i5_3_lut.init = 16'hcaca;
    LUT4 i20127_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n26823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20127_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n26867), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n26825), .SP(n2622), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i20128_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n26824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20128_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3539), .Z(n3540[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i1_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24196), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24195), .COUT(n24196), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24194), .COUT(n24195), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24193), .COUT(n24194), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24192), .COUT(n24193), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24191), .COUT(n24192), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24190), .COUT(n24191), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24189), .COUT(n24190), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24188), .COUT(n24189), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24187), .COUT(n24188), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24186), .COUT(n24187), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24185), .COUT(n24186), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24184), .COUT(n24185), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24183), .COUT(n24184), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24182), .COUT(n24183), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24181), .COUT(n24182), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n24181), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    PFUMX i20171 (.BLUT(n26865), .ALUT(n26866), .C0(\register_addr[0] ), 
          .Z(n26867));
    LUT4 i13254_2_lut (.A(Stepper_Y_Dir_c), .B(\register_addr[0] ), .Z(n7684[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13254_2_lut.init = 16'h2222;
    LUT4 mux_1755_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n5671[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1755_i6_3_lut.init = 16'hcaca;
    LUT4 i13253_2_lut (.A(Stepper_Y_En_c), .B(\register_addr[0] ), .Z(n7684[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13253_2_lut.init = 16'h2222;
    LUT4 mux_1755_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n5671[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1755_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1755_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5671[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1755_i8_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n8273), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n8273), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n8273), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n8273), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n8273), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n8273), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n8273), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n8273), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i1 (.D(n611), .SP(n13363), .CK(debug_c_c), 
            .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n12649), .CD(n11054), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n12649), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n12649), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n12649), .CD(n28477), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n12649), .PD(n28477), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n12649), .CD(n28477), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n12649), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n26540), .SP(n2622), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3540[31]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3540[30]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3540[29]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3540[28]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3540[27]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3540[26]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3540[25]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3540[24]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3540[23]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3540[22]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3540[21]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3540[20]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3540[19]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3540[18]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3540[17]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3540[16]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3540[15]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3540[14]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3540[13]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3540[12]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3540[11]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3540[10]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3540[9]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3540[8]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3540[7]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3540[6]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3540[5]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3540[4]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3540[3]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3540[2]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3540[1]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i13256_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n7684[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13256_2_lut.init = 16'h2222;
    LUT4 mux_1755_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n5671[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1755_i4_3_lut.init = 16'hcaca;
    LUT4 i20169_3_lut (.A(Stepper_Y_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n26865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20169_3_lut.init = 16'hcaca;
    LUT4 i20170_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n26866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20170_3_lut.init = 16'hcaca;
    LUT4 i20109_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n26805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20109_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1494_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3539), 
         .Z(n3540[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i32_3_lut.init = 16'hcaca;
    LUT4 i13221_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13221_4_lut.init = 16'hc088;
    LUT4 i13222_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13222_4_lut.init = 16'hc088;
    LUT4 mux_1494_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3539), 
         .Z(n3540[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i31_3_lut.init = 16'hcaca;
    LUT4 i13223_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13223_4_lut.init = 16'hc088;
    LUT4 i13224_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13224_4_lut.init = 16'hc088;
    LUT4 i13225_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13225_4_lut.init = 16'hc088;
    LUT4 i13226_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13226_4_lut.init = 16'hc088;
    LUT4 i13227_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13227_4_lut.init = 16'hc088;
    LUT4 i13228_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13228_4_lut.init = 16'hc088;
    LUT4 i13229_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13229_4_lut.init = 16'hc088;
    LUT4 i13230_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13230_4_lut.init = 16'hc088;
    LUT4 i13231_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13231_4_lut.init = 16'hc088;
    LUT4 i13232_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13232_4_lut.init = 16'hc088;
    LUT4 i13233_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13233_4_lut.init = 16'hc088;
    LUT4 mux_1494_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3539), 
         .Z(n3540[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i30_3_lut.init = 16'hcaca;
    LUT4 i13234_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13234_4_lut.init = 16'hc088;
    LUT4 mux_1494_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3539), 
         .Z(n3540[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i29_3_lut.init = 16'hcaca;
    LUT4 i13235_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13235_4_lut.init = 16'hc088;
    LUT4 mux_1494_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3539), 
         .Z(n3540[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i28_3_lut.init = 16'hcaca;
    PFUMX mux_1759_i4 (.BLUT(n7684[3]), .ALUT(n5671[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    LUT4 mux_1494_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3539), 
         .Z(n3540[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i27_3_lut.init = 16'hcaca;
    LUT4 i13236_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13236_4_lut.init = 16'hc088;
    LUT4 mux_1494_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3539), 
         .Z(n3540[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3539), 
         .Z(n3540[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i25_3_lut.init = 16'hcaca;
    LUT4 i13237_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13237_4_lut.init = 16'hc088;
    LUT4 mux_1494_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3539), 
         .Z(n3540[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3539), 
         .Z(n3540[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3539), 
         .Z(n3540[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i22_3_lut.init = 16'hcaca;
    LUT4 i13238_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13238_4_lut.init = 16'hc088;
    FD1P3AX int_step_182 (.D(n28411), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1494_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3539), 
         .Z(n3540[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3539), 
         .Z(n3540[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3539), 
         .Z(n3540[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i19_3_lut.init = 16'hcaca;
    LUT4 i13239_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13239_4_lut.init = 16'hc088;
    LUT4 i13240_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13240_4_lut.init = 16'hc088;
    LUT4 i13241_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13241_4_lut.init = 16'hc088;
    LUT4 i13242_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13242_4_lut.init = 16'hc088;
    LUT4 i13243_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13243_4_lut.init = 16'hc088;
    LUT4 i13244_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13244_4_lut.init = 16'hc088;
    LUT4 mux_1494_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3539), 
         .Z(n3540[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3539), 
         .Z(n3540[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i17_3_lut.init = 16'hcaca;
    PFUMX mux_1759_i5 (.BLUT(n7684[4]), .ALUT(n5671[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    LUT4 mux_1494_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3539), 
         .Z(n3540[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3539), 
         .Z(n3540[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3539), 
         .Z(n3540[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i14_3_lut.init = 16'hcaca;
    PFUMX mux_1759_i6 (.BLUT(n7684[5]), .ALUT(n5671[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    LUT4 mux_1494_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3539), 
         .Z(n3540[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3539), 
         .Z(n3540[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i12_3_lut.init = 16'hcaca;
    PFUMX mux_1759_i7 (.BLUT(n7684[6]), .ALUT(n5671[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    PFUMX mux_1759_i8 (.BLUT(n7685), .ALUT(n5671[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    LUT4 mux_1494_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3539), 
         .Z(n3540[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3539), .Z(n3540[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3539), .Z(n3540[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3539), .Z(n3540[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3539), .Z(n3540[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3539), .Z(n3540[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3539), .Z(n3540[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3539), .Z(n3540[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3539), .Z(n3540[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1494_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3539), .Z(n3540[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1494_i2_3_lut.init = 16'hcaca;
    LUT4 i20110_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n26806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20110_3_lut.init = 16'hcaca;
    ClockDivider_U6 step_clk_gen (.step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n28477(n28477), .div_factor_reg({div_factor_reg}), .GND_net(GND_net), 
            .n28400(n28400), .n14873(n14873), .n7244(n7244), .n7278(n7278)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U6
//

module ClockDivider_U6 (step_clk, debug_c_c, n28477, div_factor_reg, 
            GND_net, n28400, n14873, n7244, n7278) /* synthesis syn_module_defined=1 */ ;
    output step_clk;
    input debug_c_c;
    input n28477;
    input [31:0]div_factor_reg;
    input GND_net;
    input n28400;
    input n14873;
    output n7244;
    output n7278;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7209, n23922, n23923, n23921, n23920, n23919, n23918, 
        n23917, n23916, n23915, n23914, n23913, n23912;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n24344, n24343, n24342, n24341, n23911, n23910, n24340, 
        n24339, n24338, n23909, n24337, n24336, n24335, n24334, 
        n24333, n24332, n24331, n24330, n24329;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n23956, n23955, n23954, n23953, n23952, n23951, n23950, 
        n23949, n23948, n24132;
    wire [31:0]n40;
    
    wire n24131, n24130, n24129, n24128, n24127, n24126, n23947, 
        n24125, n23946, n24124, n24123, n24122, n24121, n24120, 
        n24119, n24118, n24117, n23945, n23944, n23943, n23942, 
        n23941, n23940, n23939, n23938, n23937, n23936, n23935, 
        n23934, n23933, n23932, n23931, n23930, n23929, n23928, 
        n23927, n23926, n23925, n23924;
    
    FD1S3IX clk_o_22 (.D(n7209), .CK(debug_c_c), .CD(n28477), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1874_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23922), .COUT(n23923));
    defparam sub_1874_add_2_29.INIT0 = 16'hf555;
    defparam sub_1874_add_2_29.INIT1 = 16'hf555;
    defparam sub_1874_add_2_29.INJECT1_0 = "NO";
    defparam sub_1874_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23921), .COUT(n23922));
    defparam sub_1874_add_2_27.INIT0 = 16'hf555;
    defparam sub_1874_add_2_27.INIT1 = 16'hf555;
    defparam sub_1874_add_2_27.INJECT1_0 = "NO";
    defparam sub_1874_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23920), .COUT(n23921));
    defparam sub_1874_add_2_25.INIT0 = 16'hf555;
    defparam sub_1874_add_2_25.INIT1 = 16'hf555;
    defparam sub_1874_add_2_25.INJECT1_0 = "NO";
    defparam sub_1874_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23919), .COUT(n23920));
    defparam sub_1874_add_2_23.INIT0 = 16'hf555;
    defparam sub_1874_add_2_23.INIT1 = 16'hf555;
    defparam sub_1874_add_2_23.INJECT1_0 = "NO";
    defparam sub_1874_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23918), .COUT(n23919));
    defparam sub_1874_add_2_21.INIT0 = 16'hf555;
    defparam sub_1874_add_2_21.INIT1 = 16'hf555;
    defparam sub_1874_add_2_21.INJECT1_0 = "NO";
    defparam sub_1874_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23917), .COUT(n23918));
    defparam sub_1874_add_2_19.INIT0 = 16'hf555;
    defparam sub_1874_add_2_19.INIT1 = 16'hf555;
    defparam sub_1874_add_2_19.INJECT1_0 = "NO";
    defparam sub_1874_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23916), .COUT(n23917));
    defparam sub_1874_add_2_17.INIT0 = 16'hf555;
    defparam sub_1874_add_2_17.INIT1 = 16'hf555;
    defparam sub_1874_add_2_17.INJECT1_0 = "NO";
    defparam sub_1874_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23915), .COUT(n23916));
    defparam sub_1874_add_2_15.INIT0 = 16'hf555;
    defparam sub_1874_add_2_15.INIT1 = 16'hf555;
    defparam sub_1874_add_2_15.INJECT1_0 = "NO";
    defparam sub_1874_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23914), .COUT(n23915));
    defparam sub_1874_add_2_13.INIT0 = 16'hf555;
    defparam sub_1874_add_2_13.INIT1 = 16'hf555;
    defparam sub_1874_add_2_13.INJECT1_0 = "NO";
    defparam sub_1874_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23913), .COUT(n23914));
    defparam sub_1874_add_2_11.INIT0 = 16'hf555;
    defparam sub_1874_add_2_11.INIT1 = 16'hf555;
    defparam sub_1874_add_2_11.INJECT1_0 = "NO";
    defparam sub_1874_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23912), .COUT(n23913));
    defparam sub_1874_add_2_9.INIT0 = 16'hf555;
    defparam sub_1874_add_2_9.INIT1 = 16'hf555;
    defparam sub_1874_add_2_9.INJECT1_0 = "NO";
    defparam sub_1874_add_2_9.INJECT1_1 = "NO";
    FD1S3IX count_2373__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i0.GSR = "ENABLED";
    CCU2D count_2373_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24344), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_33.INIT1 = 16'h0000;
    defparam count_2373_add_4_33.INJECT1_0 = "NO";
    defparam count_2373_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24343), .COUT(n24344), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_31.INJECT1_0 = "NO";
    defparam count_2373_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24342), .COUT(n24343), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_29.INJECT1_0 = "NO";
    defparam count_2373_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24341), .COUT(n24342), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_27.INJECT1_0 = "NO";
    defparam count_2373_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23911), .COUT(n23912));
    defparam sub_1874_add_2_7.INIT0 = 16'hf555;
    defparam sub_1874_add_2_7.INIT1 = 16'hf555;
    defparam sub_1874_add_2_7.INJECT1_0 = "NO";
    defparam sub_1874_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23910), .COUT(n23911));
    defparam sub_1874_add_2_5.INIT0 = 16'hf555;
    defparam sub_1874_add_2_5.INIT1 = 16'hf555;
    defparam sub_1874_add_2_5.INJECT1_0 = "NO";
    defparam sub_1874_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24340), .COUT(n24341), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_25.INJECT1_0 = "NO";
    defparam count_2373_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24339), .COUT(n24340), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_23.INJECT1_0 = "NO";
    defparam count_2373_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24338), .COUT(n24339), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_21.INJECT1_0 = "NO";
    defparam count_2373_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23909), .COUT(n23910));
    defparam sub_1874_add_2_3.INIT0 = 16'hf555;
    defparam sub_1874_add_2_3.INIT1 = 16'hf555;
    defparam sub_1874_add_2_3.INJECT1_0 = "NO";
    defparam sub_1874_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24337), .COUT(n24338), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_19.INJECT1_0 = "NO";
    defparam count_2373_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24336), .COUT(n24337), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_17.INJECT1_0 = "NO";
    defparam count_2373_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24335), .COUT(n24336), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_15.INJECT1_0 = "NO";
    defparam count_2373_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24334), .COUT(n24335), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_13.INJECT1_0 = "NO";
    defparam count_2373_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n23909));
    defparam sub_1874_add_2_1.INIT0 = 16'h0000;
    defparam sub_1874_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1874_add_2_1.INJECT1_0 = "NO";
    defparam sub_1874_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24333), .COUT(n24334), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_11.INJECT1_0 = "NO";
    defparam count_2373_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24332), .COUT(n24333), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_9.INJECT1_0 = "NO";
    defparam count_2373_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24331), .COUT(n24332), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_7.INJECT1_0 = "NO";
    defparam count_2373_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24330), .COUT(n24331), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_5.INJECT1_0 = "NO";
    defparam count_2373_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24329), .COUT(n24330), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2373_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2373_add_4_3.INJECT1_0 = "NO";
    defparam count_2373_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2373_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24329), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373_add_4_1.INIT0 = 16'hF000;
    defparam count_2373_add_4_1.INIT1 = 16'h0555;
    defparam count_2373_add_4_1.INJECT1_0 = "NO";
    defparam count_2373_add_4_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    CCU2D sub_1871_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23956), .S1(n7209));
    defparam sub_1871_add_2_33.INIT0 = 16'h5555;
    defparam sub_1871_add_2_33.INIT1 = 16'h0000;
    defparam sub_1871_add_2_33.INJECT1_0 = "NO";
    defparam sub_1871_add_2_33.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28400), .PD(n14873), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_1871_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23955), .COUT(n23956));
    defparam sub_1871_add_2_31.INIT0 = 16'h5999;
    defparam sub_1871_add_2_31.INIT1 = 16'h5999;
    defparam sub_1871_add_2_31.INJECT1_0 = "NO";
    defparam sub_1871_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23954), .COUT(n23955));
    defparam sub_1871_add_2_29.INIT0 = 16'h5999;
    defparam sub_1871_add_2_29.INIT1 = 16'h5999;
    defparam sub_1871_add_2_29.INJECT1_0 = "NO";
    defparam sub_1871_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23953), .COUT(n23954));
    defparam sub_1871_add_2_27.INIT0 = 16'h5999;
    defparam sub_1871_add_2_27.INIT1 = 16'h5999;
    defparam sub_1871_add_2_27.INJECT1_0 = "NO";
    defparam sub_1871_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23952), .COUT(n23953));
    defparam sub_1871_add_2_25.INIT0 = 16'h5999;
    defparam sub_1871_add_2_25.INIT1 = 16'h5999;
    defparam sub_1871_add_2_25.INJECT1_0 = "NO";
    defparam sub_1871_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23951), .COUT(n23952));
    defparam sub_1871_add_2_23.INIT0 = 16'h5999;
    defparam sub_1871_add_2_23.INIT1 = 16'h5999;
    defparam sub_1871_add_2_23.INJECT1_0 = "NO";
    defparam sub_1871_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23950), .COUT(n23951));
    defparam sub_1871_add_2_21.INIT0 = 16'h5999;
    defparam sub_1871_add_2_21.INIT1 = 16'h5999;
    defparam sub_1871_add_2_21.INJECT1_0 = "NO";
    defparam sub_1871_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23949), .COUT(n23950));
    defparam sub_1871_add_2_19.INIT0 = 16'h5999;
    defparam sub_1871_add_2_19.INIT1 = 16'h5999;
    defparam sub_1871_add_2_19.INJECT1_0 = "NO";
    defparam sub_1871_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23948), .COUT(n23949));
    defparam sub_1871_add_2_17.INIT0 = 16'h5999;
    defparam sub_1871_add_2_17.INIT1 = 16'h5999;
    defparam sub_1871_add_2_17.INJECT1_0 = "NO";
    defparam sub_1871_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24132), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24131), .COUT(n24132), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24130), .COUT(n24131), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24129), .COUT(n24130), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24128), .COUT(n24129), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24127), .COUT(n24128), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24126), .COUT(n24127), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23947), .COUT(n23948));
    defparam sub_1871_add_2_15.INIT0 = 16'h5999;
    defparam sub_1871_add_2_15.INIT1 = 16'h5999;
    defparam sub_1871_add_2_15.INJECT1_0 = "NO";
    defparam sub_1871_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24125), .COUT(n24126), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23946), .COUT(n23947));
    defparam sub_1871_add_2_13.INIT0 = 16'h5999;
    defparam sub_1871_add_2_13.INIT1 = 16'h5999;
    defparam sub_1871_add_2_13.INJECT1_0 = "NO";
    defparam sub_1871_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24124), .COUT(n24125), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24123), .COUT(n24124), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24122), .COUT(n24123), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24121), .COUT(n24122), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24120), .COUT(n24121), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24119), .COUT(n24120), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24118), .COUT(n24119), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24117), .COUT(n24118), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23945), .COUT(n23946));
    defparam sub_1871_add_2_11.INIT0 = 16'h5999;
    defparam sub_1871_add_2_11.INIT1 = 16'h5999;
    defparam sub_1871_add_2_11.INJECT1_0 = "NO";
    defparam sub_1871_add_2_11.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28400), .CD(n14873), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_1871_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23944), .COUT(n23945));
    defparam sub_1871_add_2_9.INIT0 = 16'h5999;
    defparam sub_1871_add_2_9.INIT1 = 16'h5999;
    defparam sub_1871_add_2_9.INJECT1_0 = "NO";
    defparam sub_1871_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23943), .COUT(n23944));
    defparam sub_1871_add_2_7.INIT0 = 16'h5999;
    defparam sub_1871_add_2_7.INIT1 = 16'h5999;
    defparam sub_1871_add_2_7.INJECT1_0 = "NO";
    defparam sub_1871_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24117), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23942), .COUT(n23943));
    defparam sub_1871_add_2_5.INIT0 = 16'h5999;
    defparam sub_1871_add_2_5.INIT1 = 16'h5999;
    defparam sub_1871_add_2_5.INJECT1_0 = "NO";
    defparam sub_1871_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1871_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23941), .COUT(n23942));
    defparam sub_1871_add_2_3.INIT0 = 16'h5999;
    defparam sub_1871_add_2_3.INIT1 = 16'h5999;
    defparam sub_1871_add_2_3.INJECT1_0 = "NO";
    defparam sub_1871_add_2_3.INJECT1_1 = "NO";
    FD1S3IX count_2373__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i1.GSR = "ENABLED";
    CCU2D sub_1871_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n23941));
    defparam sub_1871_add_2_1.INIT0 = 16'h0000;
    defparam sub_1871_add_2_1.INIT1 = 16'h5999;
    defparam sub_1871_add_2_1.INJECT1_0 = "NO";
    defparam sub_1871_add_2_1.INJECT1_1 = "NO";
    FD1S3IX count_2373__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i2.GSR = "ENABLED";
    FD1S3IX count_2373__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i3.GSR = "ENABLED";
    FD1S3IX count_2373__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i4.GSR = "ENABLED";
    FD1S3IX count_2373__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i5.GSR = "ENABLED";
    FD1S3IX count_2373__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i6.GSR = "ENABLED";
    FD1S3IX count_2373__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i7.GSR = "ENABLED";
    FD1S3IX count_2373__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i8.GSR = "ENABLED";
    FD1S3IX count_2373__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i9.GSR = "ENABLED";
    FD1S3IX count_2373__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i10.GSR = "ENABLED";
    FD1S3IX count_2373__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i11.GSR = "ENABLED";
    FD1S3IX count_2373__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i12.GSR = "ENABLED";
    FD1S3IX count_2373__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i13.GSR = "ENABLED";
    FD1S3IX count_2373__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i14.GSR = "ENABLED";
    FD1S3IX count_2373__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i15.GSR = "ENABLED";
    FD1S3IX count_2373__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i16.GSR = "ENABLED";
    FD1S3IX count_2373__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i17.GSR = "ENABLED";
    FD1S3IX count_2373__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i18.GSR = "ENABLED";
    FD1S3IX count_2373__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i19.GSR = "ENABLED";
    FD1S3IX count_2373__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i20.GSR = "ENABLED";
    FD1S3IX count_2373__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i21.GSR = "ENABLED";
    FD1S3IX count_2373__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i22.GSR = "ENABLED";
    FD1S3IX count_2373__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i23.GSR = "ENABLED";
    FD1S3IX count_2373__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i24.GSR = "ENABLED";
    FD1S3IX count_2373__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i25.GSR = "ENABLED";
    FD1S3IX count_2373__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i26.GSR = "ENABLED";
    FD1S3IX count_2373__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i27.GSR = "ENABLED";
    FD1S3IX count_2373__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i28.GSR = "ENABLED";
    FD1S3IX count_2373__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i29.GSR = "ENABLED";
    FD1S3IX count_2373__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i30.GSR = "ENABLED";
    FD1S3IX count_2373__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28400), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2373__i31.GSR = "ENABLED";
    CCU2D sub_1873_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23940), .S1(n7244));
    defparam sub_1873_add_2_33.INIT0 = 16'h5999;
    defparam sub_1873_add_2_33.INIT1 = 16'h0000;
    defparam sub_1873_add_2_33.INJECT1_0 = "NO";
    defparam sub_1873_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23939), .COUT(n23940));
    defparam sub_1873_add_2_31.INIT0 = 16'h5999;
    defparam sub_1873_add_2_31.INIT1 = 16'h5999;
    defparam sub_1873_add_2_31.INJECT1_0 = "NO";
    defparam sub_1873_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23938), .COUT(n23939));
    defparam sub_1873_add_2_29.INIT0 = 16'h5999;
    defparam sub_1873_add_2_29.INIT1 = 16'h5999;
    defparam sub_1873_add_2_29.INJECT1_0 = "NO";
    defparam sub_1873_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23937), .COUT(n23938));
    defparam sub_1873_add_2_27.INIT0 = 16'h5999;
    defparam sub_1873_add_2_27.INIT1 = 16'h5999;
    defparam sub_1873_add_2_27.INJECT1_0 = "NO";
    defparam sub_1873_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23936), .COUT(n23937));
    defparam sub_1873_add_2_25.INIT0 = 16'h5999;
    defparam sub_1873_add_2_25.INIT1 = 16'h5999;
    defparam sub_1873_add_2_25.INJECT1_0 = "NO";
    defparam sub_1873_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23935), .COUT(n23936));
    defparam sub_1873_add_2_23.INIT0 = 16'h5999;
    defparam sub_1873_add_2_23.INIT1 = 16'h5999;
    defparam sub_1873_add_2_23.INJECT1_0 = "NO";
    defparam sub_1873_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23934), .COUT(n23935));
    defparam sub_1873_add_2_21.INIT0 = 16'h5999;
    defparam sub_1873_add_2_21.INIT1 = 16'h5999;
    defparam sub_1873_add_2_21.INJECT1_0 = "NO";
    defparam sub_1873_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23933), .COUT(n23934));
    defparam sub_1873_add_2_19.INIT0 = 16'h5999;
    defparam sub_1873_add_2_19.INIT1 = 16'h5999;
    defparam sub_1873_add_2_19.INJECT1_0 = "NO";
    defparam sub_1873_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23932), .COUT(n23933));
    defparam sub_1873_add_2_17.INIT0 = 16'h5999;
    defparam sub_1873_add_2_17.INIT1 = 16'h5999;
    defparam sub_1873_add_2_17.INJECT1_0 = "NO";
    defparam sub_1873_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23931), .COUT(n23932));
    defparam sub_1873_add_2_15.INIT0 = 16'h5999;
    defparam sub_1873_add_2_15.INIT1 = 16'h5999;
    defparam sub_1873_add_2_15.INJECT1_0 = "NO";
    defparam sub_1873_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23930), .COUT(n23931));
    defparam sub_1873_add_2_13.INIT0 = 16'h5999;
    defparam sub_1873_add_2_13.INIT1 = 16'h5999;
    defparam sub_1873_add_2_13.INJECT1_0 = "NO";
    defparam sub_1873_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23929), .COUT(n23930));
    defparam sub_1873_add_2_11.INIT0 = 16'h5999;
    defparam sub_1873_add_2_11.INIT1 = 16'h5999;
    defparam sub_1873_add_2_11.INJECT1_0 = "NO";
    defparam sub_1873_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23928), .COUT(n23929));
    defparam sub_1873_add_2_9.INIT0 = 16'h5999;
    defparam sub_1873_add_2_9.INIT1 = 16'h5999;
    defparam sub_1873_add_2_9.INJECT1_0 = "NO";
    defparam sub_1873_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23927), .COUT(n23928));
    defparam sub_1873_add_2_7.INIT0 = 16'h5999;
    defparam sub_1873_add_2_7.INIT1 = 16'h5999;
    defparam sub_1873_add_2_7.INJECT1_0 = "NO";
    defparam sub_1873_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23926), .COUT(n23927));
    defparam sub_1873_add_2_5.INIT0 = 16'h5999;
    defparam sub_1873_add_2_5.INIT1 = 16'h5999;
    defparam sub_1873_add_2_5.INJECT1_0 = "NO";
    defparam sub_1873_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23925), .COUT(n23926));
    defparam sub_1873_add_2_3.INIT0 = 16'h5999;
    defparam sub_1873_add_2_3.INIT1 = 16'h5999;
    defparam sub_1873_add_2_3.INJECT1_0 = "NO";
    defparam sub_1873_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1873_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n23925));
    defparam sub_1873_add_2_1.INIT0 = 16'h0000;
    defparam sub_1873_add_2_1.INIT1 = 16'h5999;
    defparam sub_1873_add_2_1.INJECT1_0 = "NO";
    defparam sub_1873_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23924), .S1(n7278));
    defparam sub_1874_add_2_33.INIT0 = 16'hf555;
    defparam sub_1874_add_2_33.INIT1 = 16'h0000;
    defparam sub_1874_add_2_33.INJECT1_0 = "NO";
    defparam sub_1874_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1874_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23923), .COUT(n23924));
    defparam sub_1874_add_2_31.INIT0 = 16'hf555;
    defparam sub_1874_add_2_31.INIT1 = 16'hf555;
    defparam sub_1874_add_2_31.INJECT1_0 = "NO";
    defparam sub_1874_add_2_31.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (\register_addr[1] , \register_addr[0] , 
            read_value, debug_c_c, n12599, GND_net, n28477, databus, 
            n3356, n32, prev_step_clk, step_clk, n22, VCC_net, Stepper_A_nFault_c, 
            \read_size[0] , n26437, Stepper_A_M0_c_0, n12795, n579, 
            limit_latched, prev_limit_latched, n12781, prev_select, 
            n28476, n28441, n608, n610, \control_reg[7] , n28442, 
            n10107, Stepper_A_En_c, Stepper_A_Dir_c, Stepper_A_M2_c_2, 
            Stepper_A_M1_c_1, \read_size[2] , n26439, n32_adj_1, prev_step_clk_adj_2, 
            step_clk_adj_3, n28410, n22_adj_4, n28411, n32_adj_5, 
            limit_c_3, n24744, Stepper_A_Step_c, n7703, n28399, n14876, 
            n7486, n7452) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[1] ;
    input \register_addr[0] ;
    output [31:0]read_value;
    input debug_c_c;
    input n12599;
    input GND_net;
    input n28477;
    input [31:0]databus;
    input n3356;
    input n32;
    input prev_step_clk;
    input step_clk;
    output n22;
    input VCC_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n26437;
    output Stepper_A_M0_c_0;
    input n12795;
    input n579;
    output limit_latched;
    output prev_limit_latched;
    input n12781;
    output prev_select;
    input n28476;
    input n28441;
    input n608;
    input n610;
    output \control_reg[7] ;
    input n28442;
    input n10107;
    output Stepper_A_En_c;
    output Stepper_A_Dir_c;
    output Stepper_A_M2_c_2;
    output Stepper_A_M1_c_1;
    output \read_size[2] ;
    input n26439;
    input n32_adj_1;
    input prev_step_clk_adj_2;
    input step_clk_adj_3;
    output n28410;
    output n22_adj_4;
    output n28411;
    input n32_adj_5;
    input limit_c_3;
    output n24744;
    output Stepper_A_Step_c;
    input n7703;
    input n28399;
    input n14876;
    output n7486;
    output n7452;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n11;
    wire [31:0]n100;
    
    wire n26811, n26812, n26813, n26814, n26815, n26816;
    wire [31:0]n99;
    wire [31:0]n3357;
    wire [31:0]n224;
    
    wire fault_latched, prev_step_clk_adj_15, step_clk_adj_16, n182;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n26861, n26859, n26860, n24164, n24163, n24162, n24161, 
        n24160, n24159, n24158, n24157, n24156, n24155, n24154, 
        n24153;
    wire [7:0]n7702;
    
    wire n24152;
    wire [31:0]n6299;
    
    wire n24151, n24150, n24149, n49_adj_22, n62_adj_23, n58_adj_24, 
        n50, n41_adj_25, n60_adj_26, n54_adj_27, n42, n52, n38, 
        n56, n46, n28413, n22_adj_28, int_step;
    
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[20]), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n11)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i13199_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13199_4_lut.init = 16'hc088;
    LUT4 i13200_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13200_4_lut.init = 16'hc088;
    LUT4 i13201_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13201_4_lut.init = 16'hc088;
    PFUMX i20117 (.BLUT(n26811), .ALUT(n26812), .C0(\register_addr[1] ), 
          .Z(n26813));
    LUT4 i13202_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13202_4_lut.init = 16'hc088;
    LUT4 i13203_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13203_4_lut.init = 16'hc088;
    PFUMX i20120 (.BLUT(n26814), .ALUT(n26815), .C0(\register_addr[0] ), 
          .Z(n26816));
    LUT4 i13204_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13204_4_lut.init = 16'hc088;
    FD1P3IX read_value__i0 (.D(n26813), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i13205_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13205_4_lut.init = 16'hc088;
    LUT4 i13206_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13206_4_lut.init = 16'hc088;
    LUT4 i13207_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13207_4_lut.init = 16'hc088;
    LUT4 i13208_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13208_4_lut.init = 16'hc088;
    LUT4 i13209_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13209_4_lut.init = 16'hc088;
    LUT4 i13210_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13210_4_lut.init = 16'hc088;
    LUT4 i13617_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n99[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13617_4_lut.init = 16'hc088;
    LUT4 i13610_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n99[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13610_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_2 (.A(\register_addr[1] ), .B(div_factor_reg[24]), 
         .C(steps_reg[24]), .D(\register_addr[0] ), .Z(n99[24])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_2.init = 16'ha088;
    LUT4 i13609_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n99[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13609_4_lut.init = 16'hc088;
    LUT4 i13608_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n99[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13608_4_lut.init = 16'hc088;
    FD1S3IX steps_reg__i25 (.D(n3357[25]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    LUT4 i13607_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n99[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13607_4_lut.init = 16'hc088;
    LUT4 i13606_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n99[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13606_4_lut.init = 16'hc088;
    LUT4 i13605_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n99[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13605_4_lut.init = 16'hc088;
    LUT4 i13604_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n99[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13604_4_lut.init = 16'hc088;
    FD1S3IX steps_reg__i24 (.D(n3357[24]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    LUT4 i13603_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n99[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i13603_4_lut.init = 16'hc088;
    FD1S3IX steps_reg__i23 (.D(n3357[23]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3357[22]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3357[21]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3357[20]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3357[19]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3357[18]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3357[17]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3357[16]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    LUT4 mux_1447_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3356), 
         .Z(n3357[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3356), 
         .Z(n3357[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i23_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i15 (.D(n3357[15]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3357[14]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3357[0]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut (.A(n32), .B(prev_step_clk), .C(step_clk), .D(n28477), 
         .Z(n22)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut.init = 16'h002c;
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3357[13]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3357[12]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    LUT4 mux_1447_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3356), 
         .Z(n3357[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i22_3_lut.init = 16'hcaca;
    FD1P3AX read_size__i1 (.D(n26437), .SP(n12599), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12795), .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk_adj_16), .CK(debug_c_c), .Q(prev_step_clk_adj_15)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12781), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3357[11]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n28476), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3357[10]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3357[9]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3357[8]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3357[7]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3357[6]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3357[5]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3357[4]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3357[3]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3357[2]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3357[1]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1447_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3356), 
         .Z(n3357[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3356), 
         .Z(n3357[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3356), 
         .Z(n3357[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i19_3_lut.init = 16'hcaca;
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n28441), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n28441), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n28441), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n28441), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n28441), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n28441), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n28441), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n12781), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12781), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n28442), .CD(n10107), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n28442), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n28442), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n12795), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n28442), .PD(n28477), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n12795), .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n28442), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n26439), .SP(n12599), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3357[31]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3357[30]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3357[29]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3357[28]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3357[27]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3357[26]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n11), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n12599), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n26861), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n26816), .SP(n12599), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_289 (.A(n32_adj_1), .B(prev_step_clk_adj_2), .C(step_clk_adj_3), 
         .Z(n28410)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_289.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_adj_3 (.A(n32_adj_1), .B(prev_step_clk_adj_2), .C(step_clk_adj_3), 
         .D(n28477), .Z(n22_adj_4)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_3.init = 16'h002c;
    LUT4 i2_3_lut_rep_290 (.A(n32), .B(prev_step_clk), .C(step_clk), .Z(n28411)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_290.init = 16'h2020;
    LUT4 mux_1447_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3356), 
         .Z(n3357[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3356), 
         .Z(n3357[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i17_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    LUT4 mux_1447_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3356), 
         .Z(n3357[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i26_3_lut.init = 16'hcaca;
    PFUMX i20165 (.BLUT(n26859), .ALUT(n26860), .C0(\register_addr[0] ), 
          .Z(n26861));
    LUT4 mux_1447_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3356), 
         .Z(n3357[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3356), 
         .Z(n3357[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3356), 
         .Z(n3357[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3356), .Z(n3357[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i1_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24164), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24163), .COUT(n24164), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24162), .COUT(n24163), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24161), .COUT(n24162), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24160), .COUT(n24161), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24159), .COUT(n24160), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24158), .COUT(n24159), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24157), .COUT(n24158), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24156), .COUT(n24157), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24155), .COUT(n24156), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24154), .COUT(n24155), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24153), .COUT(n24154), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    LUT4 i13197_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n7702[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13197_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24152), .COUT(n24153), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 mux_1807_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n6299[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1807_i4_3_lut.init = 16'hcaca;
    LUT4 i13196_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7702[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13196_2_lut.init = 16'h2222;
    LUT4 i12261_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n6299[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i12261_3_lut.init = 16'hcaca;
    LUT4 i13195_2_lut (.A(Stepper_A_Dir_c), .B(\register_addr[0] ), .Z(n7702[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13195_2_lut.init = 16'h2222;
    LUT4 mux_1807_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n6299[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1807_i6_3_lut.init = 16'hcaca;
    LUT4 i13194_2_lut (.A(Stepper_A_En_c), .B(\register_addr[0] ), .Z(n7702[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13194_2_lut.init = 16'h2222;
    LUT4 mux_1807_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n6299[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1807_i7_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    LUT4 mux_1807_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6299[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1807_i8_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24151), .COUT(n24152), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    LUT4 mux_1447_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3356), 
         .Z(n3357[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3356), 
         .Z(n3357[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i13_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24150), .COUT(n24151), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24149), .COUT(n24150), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32_adj_5), .C1(step_clk_adj_16), .D1(prev_step_clk_adj_15), 
          .COUT(n24149), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i20118_3_lut (.A(Stepper_A_M1_c_1), .B(div_factor_reg[1]), .C(\register_addr[1] ), 
         .Z(n26814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20118_3_lut.init = 16'hcaca;
    LUT4 i13198_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13198_4_lut.init = 16'hc088;
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i20163_3_lut (.A(Stepper_A_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n26859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20163_3_lut.init = 16'hcaca;
    LUT4 i20164_3_lut (.A(n32_adj_5), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n26860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20164_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49_adj_22), .B(n62_adj_23), .C(n58_adj_24), .D(n50), 
         .Z(n24744)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[20]), .Z(n49_adj_22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41_adj_25), .B(n60_adj_26), .C(n54_adj_27), .D(n42), 
         .Z(n62_adj_23)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[8]), 
         .Z(n58_adj_24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[4]), .B(steps_reg[0]), .Z(n41_adj_25)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[22]), .B(n56), .C(n46), .D(steps_reg[9]), 
         .Z(n60_adj_26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[26]), .B(steps_reg[1]), .C(steps_reg[29]), 
         .D(steps_reg[18]), .Z(n54_adj_27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[2]), .B(steps_reg[25]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[5]), .B(steps_reg[10]), .C(steps_reg[6]), 
         .D(steps_reg[3]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 mux_1447_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3356), 
         .Z(n3357[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i12_3_lut.init = 16'hcaca;
    LUT4 i14_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 mux_1447_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3356), 
         .Z(n3357[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i11_3_lut.init = 16'hcaca;
    LUT4 i20_4_lut (.A(steps_reg[28]), .B(steps_reg[7]), .C(steps_reg[30]), 
         .D(steps_reg[24]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[16]), .B(steps_reg[13]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1447_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3356), .Z(n3357[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i10_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    LUT4 mux_1447_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3356), .Z(n3357[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3356), .Z(n3357[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3356), .Z(n3357[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3356), .Z(n3357[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3356), .Z(n3357[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3356), .Z(n3357[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i4_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    LUT4 mux_1447_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3356), .Z(n3357[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3356), .Z(n3357[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i2_3_lut.init = 16'hcaca;
    LUT4 i20119_3_lut (.A(fault_latched), .B(steps_reg[1]), .C(\register_addr[1] ), 
         .Z(n26815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20119_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_292 (.A(n32_adj_5), .B(prev_step_clk_adj_15), .C(step_clk_adj_16), 
         .Z(n28413)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_292.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_adj_4 (.A(n32_adj_5), .B(prev_step_clk_adj_15), 
         .C(step_clk_adj_16), .D(n28477), .Z(n22_adj_28)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_4.init = 16'h002c;
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12781), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    FD1P3AX read_value__i22 (.D(n99[22]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n99[23]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n99[24]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n99[25]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n99[26]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n99[27]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n99[28]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n99[29]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n99[30]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n99[31]), .SP(n12599), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n28413), .SP(n22_adj_28), .CK(debug_c_c), 
            .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1447_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3356), 
         .Z(n3357[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i32_3_lut.init = 16'hcaca;
    PFUMX mux_1811_i4 (.BLUT(n7702[3]), .ALUT(n6299[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_1811_i5 (.BLUT(n7702[4]), .ALUT(n6299[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1811_i6 (.BLUT(n7702[5]), .ALUT(n6299[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1811_i7 (.BLUT(n7702[6]), .ALUT(n6299[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    LUT4 mux_1447_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3356), 
         .Z(n3357[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3356), 
         .Z(n3357[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3356), 
         .Z(n3357[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1447_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3356), 
         .Z(n3357[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i28_3_lut.init = 16'hcaca;
    PFUMX mux_1811_i8 (.BLUT(n7703), .ALUT(n6299[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    LUT4 mux_1447_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3356), 
         .Z(n3357[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1447_i27_3_lut.init = 16'hcaca;
    LUT4 i20115_3_lut (.A(Stepper_A_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n26811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20115_3_lut.init = 16'hcaca;
    LUT4 i20116_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n26812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20116_3_lut.init = 16'hcaca;
    ClockDivider_U8 step_clk_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .n28399(n28399), .n14876(n14876), .div_factor_reg({div_factor_reg}), 
            .step_clk(step_clk_adj_16), .n28477(n28477), .n7486(n7486), 
            .n7452(n7452)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (GND_net, debug_c_c, n28399, n14876, div_factor_reg, 
            step_clk, n28477, n7486, n7452) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n28399;
    input n14876;
    input [31:0]div_factor_reg;
    output step_clk;
    input n28477;
    output n7486;
    output n7452;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n23825;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n40;
    
    wire n23826, n23815, n23816, n23824, n23844, n7417, n23814, 
        n23843;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n23813, n23823, n23842, n23841, n23840, n23839, n23838;
    wire [31:0]n134;
    
    wire n23837, n23836, n23822, n23835, n23821, n23834, n23833, 
        n23818, n23819, n24280, n24279, n24278, n24277, n23832, 
        n24276, n23820, n23831, n24275, n24274, n24273, n23830, 
        n24272, n24271, n24270, n24269, n24268, n24267, n23829, 
        n24266, n24265, n23817, n24100, n24099, n24098, n24097, 
        n24440, n24096, n24439, n24095, n24438, n24437, n24436, 
        n24094, n24435, n24093, n24092, n24434, n24091, n24090, 
        n24433, n24432, n24431, n24089, n24088, n24430, n24429, 
        n24087, n24428, n24427, n24426, n24086, n24425, n24085, 
        n23828, n23827;
    
    CCU2D sub_1883_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23825), .COUT(n23826));
    defparam sub_1883_add_2_27.INIT0 = 16'h5999;
    defparam sub_1883_add_2_27.INIT1 = 16'h5999;
    defparam sub_1883_add_2_27.INJECT1_0 = "NO";
    defparam sub_1883_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23815), .COUT(n23816));
    defparam sub_1883_add_2_7.INIT0 = 16'h5999;
    defparam sub_1883_add_2_7.INIT1 = 16'h5999;
    defparam sub_1883_add_2_7.INJECT1_0 = "NO";
    defparam sub_1883_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23824), .COUT(n23825));
    defparam sub_1883_add_2_25.INIT0 = 16'h5999;
    defparam sub_1883_add_2_25.INIT1 = 16'h5999;
    defparam sub_1883_add_2_25.INJECT1_0 = "NO";
    defparam sub_1883_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23844), .S1(n7417));
    defparam sub_1881_add_2_33.INIT0 = 16'h5555;
    defparam sub_1881_add_2_33.INIT1 = 16'h0000;
    defparam sub_1881_add_2_33.INJECT1_0 = "NO";
    defparam sub_1881_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23814), .COUT(n23815));
    defparam sub_1883_add_2_5.INIT0 = 16'h5999;
    defparam sub_1883_add_2_5.INIT1 = 16'h5999;
    defparam sub_1883_add_2_5.INJECT1_0 = "NO";
    defparam sub_1883_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23843), .COUT(n23844));
    defparam sub_1881_add_2_31.INIT0 = 16'h5999;
    defparam sub_1881_add_2_31.INIT1 = 16'h5999;
    defparam sub_1881_add_2_31.INJECT1_0 = "NO";
    defparam sub_1881_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23813), .COUT(n23814));
    defparam sub_1883_add_2_3.INIT0 = 16'h5999;
    defparam sub_1883_add_2_3.INIT1 = 16'h5999;
    defparam sub_1883_add_2_3.INJECT1_0 = "NO";
    defparam sub_1883_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n23813));
    defparam sub_1883_add_2_1.INIT0 = 16'h0000;
    defparam sub_1883_add_2_1.INIT1 = 16'h5999;
    defparam sub_1883_add_2_1.INJECT1_0 = "NO";
    defparam sub_1883_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23823), .COUT(n23824));
    defparam sub_1883_add_2_23.INIT0 = 16'h5999;
    defparam sub_1883_add_2_23.INIT1 = 16'h5999;
    defparam sub_1883_add_2_23.INJECT1_0 = "NO";
    defparam sub_1883_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23842), .COUT(n23843));
    defparam sub_1881_add_2_29.INIT0 = 16'h5999;
    defparam sub_1881_add_2_29.INIT1 = 16'h5999;
    defparam sub_1881_add_2_29.INJECT1_0 = "NO";
    defparam sub_1881_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23841), .COUT(n23842));
    defparam sub_1881_add_2_27.INIT0 = 16'h5999;
    defparam sub_1881_add_2_27.INIT1 = 16'h5999;
    defparam sub_1881_add_2_27.INJECT1_0 = "NO";
    defparam sub_1881_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23840), .COUT(n23841));
    defparam sub_1881_add_2_25.INIT0 = 16'h5999;
    defparam sub_1881_add_2_25.INIT1 = 16'h5999;
    defparam sub_1881_add_2_25.INJECT1_0 = "NO";
    defparam sub_1881_add_2_25.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    CCU2D sub_1881_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23839), .COUT(n23840));
    defparam sub_1881_add_2_23.INIT0 = 16'h5999;
    defparam sub_1881_add_2_23.INIT1 = 16'h5999;
    defparam sub_1881_add_2_23.INJECT1_0 = "NO";
    defparam sub_1881_add_2_23.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1S3IX clk_o_22 (.D(n7417), .CK(debug_c_c), .CD(n28477), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    CCU2D sub_1881_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23838), .COUT(n23839));
    defparam sub_1881_add_2_21.INIT0 = 16'h5999;
    defparam sub_1881_add_2_21.INIT1 = 16'h5999;
    defparam sub_1881_add_2_21.INJECT1_0 = "NO";
    defparam sub_1881_add_2_21.INJECT1_1 = "NO";
    FD1S3IX count_2375__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i0.GSR = "ENABLED";
    CCU2D sub_1881_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23837), .COUT(n23838));
    defparam sub_1881_add_2_19.INIT0 = 16'h5999;
    defparam sub_1881_add_2_19.INIT1 = 16'h5999;
    defparam sub_1881_add_2_19.INJECT1_0 = "NO";
    defparam sub_1881_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23836), .COUT(n23837));
    defparam sub_1881_add_2_17.INIT0 = 16'h5999;
    defparam sub_1881_add_2_17.INIT1 = 16'h5999;
    defparam sub_1881_add_2_17.INJECT1_0 = "NO";
    defparam sub_1881_add_2_17.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28399), .PD(n14876), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_1883_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23822), .COUT(n23823));
    defparam sub_1883_add_2_21.INIT0 = 16'h5999;
    defparam sub_1883_add_2_21.INIT1 = 16'h5999;
    defparam sub_1883_add_2_21.INJECT1_0 = "NO";
    defparam sub_1883_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23835), .COUT(n23836));
    defparam sub_1881_add_2_15.INIT0 = 16'h5999;
    defparam sub_1881_add_2_15.INIT1 = 16'h5999;
    defparam sub_1881_add_2_15.INJECT1_0 = "NO";
    defparam sub_1881_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23821), .COUT(n23822));
    defparam sub_1883_add_2_19.INIT0 = 16'h5999;
    defparam sub_1883_add_2_19.INIT1 = 16'h5999;
    defparam sub_1883_add_2_19.INJECT1_0 = "NO";
    defparam sub_1883_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23834), .COUT(n23835));
    defparam sub_1881_add_2_13.INIT0 = 16'h5999;
    defparam sub_1881_add_2_13.INIT1 = 16'h5999;
    defparam sub_1881_add_2_13.INJECT1_0 = "NO";
    defparam sub_1881_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23833), .COUT(n23834));
    defparam sub_1881_add_2_11.INIT0 = 16'h5999;
    defparam sub_1881_add_2_11.INIT1 = 16'h5999;
    defparam sub_1881_add_2_11.INJECT1_0 = "NO";
    defparam sub_1881_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23818), .COUT(n23819));
    defparam sub_1883_add_2_13.INIT0 = 16'h5999;
    defparam sub_1883_add_2_13.INIT1 = 16'h5999;
    defparam sub_1883_add_2_13.INJECT1_0 = "NO";
    defparam sub_1883_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24280), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_33.INIT1 = 16'h0000;
    defparam count_2375_add_4_33.INJECT1_0 = "NO";
    defparam count_2375_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24279), .COUT(n24280), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_31.INJECT1_0 = "NO";
    defparam count_2375_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24278), .COUT(n24279), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_29.INJECT1_0 = "NO";
    defparam count_2375_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24277), .COUT(n24278), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_27.INJECT1_0 = "NO";
    defparam count_2375_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23832), .COUT(n23833));
    defparam sub_1881_add_2_9.INIT0 = 16'h5999;
    defparam sub_1881_add_2_9.INIT1 = 16'h5999;
    defparam sub_1881_add_2_9.INJECT1_0 = "NO";
    defparam sub_1881_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24276), .COUT(n24277), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_25.INJECT1_0 = "NO";
    defparam count_2375_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23820), .COUT(n23821));
    defparam sub_1883_add_2_17.INIT0 = 16'h5999;
    defparam sub_1883_add_2_17.INIT1 = 16'h5999;
    defparam sub_1883_add_2_17.INJECT1_0 = "NO";
    defparam sub_1883_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23831), .COUT(n23832));
    defparam sub_1881_add_2_7.INIT0 = 16'h5999;
    defparam sub_1881_add_2_7.INIT1 = 16'h5999;
    defparam sub_1881_add_2_7.INJECT1_0 = "NO";
    defparam sub_1881_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24275), .COUT(n24276), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_23.INJECT1_0 = "NO";
    defparam count_2375_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24274), .COUT(n24275), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_21.INJECT1_0 = "NO";
    defparam count_2375_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24273), .COUT(n24274), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_19.INJECT1_0 = "NO";
    defparam count_2375_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23830), .COUT(n23831));
    defparam sub_1881_add_2_5.INIT0 = 16'h5999;
    defparam sub_1881_add_2_5.INIT1 = 16'h5999;
    defparam sub_1881_add_2_5.INJECT1_0 = "NO";
    defparam sub_1881_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24272), .COUT(n24273), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_17.INJECT1_0 = "NO";
    defparam count_2375_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24271), .COUT(n24272), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_15.INJECT1_0 = "NO";
    defparam count_2375_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24270), .COUT(n24271), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_13.INJECT1_0 = "NO";
    defparam count_2375_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24269), .COUT(n24270), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_11.INJECT1_0 = "NO";
    defparam count_2375_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24268), .COUT(n24269), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_9.INJECT1_0 = "NO";
    defparam count_2375_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24267), .COUT(n24268), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_7.INJECT1_0 = "NO";
    defparam count_2375_add_4_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28399), .CD(n14876), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_1881_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23829), .COUT(n23830));
    defparam sub_1881_add_2_3.INIT0 = 16'h5999;
    defparam sub_1881_add_2_3.INIT1 = 16'h5999;
    defparam sub_1881_add_2_3.INJECT1_0 = "NO";
    defparam sub_1881_add_2_3.INJECT1_1 = "NO";
    FD1S3IX count_2375__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i1.GSR = "ENABLED";
    CCU2D count_2375_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24266), .COUT(n24267), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_5.INJECT1_0 = "NO";
    defparam count_2375_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24265), .COUT(n24266), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2375_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2375_add_4_3.INJECT1_0 = "NO";
    defparam count_2375_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2375_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24265), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375_add_4_1.INIT0 = 16'hF000;
    defparam count_2375_add_4_1.INIT1 = 16'h0555;
    defparam count_2375_add_4_1.INJECT1_0 = "NO";
    defparam count_2375_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2375__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i2.GSR = "ENABLED";
    FD1S3IX count_2375__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i3.GSR = "ENABLED";
    FD1S3IX count_2375__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i4.GSR = "ENABLED";
    FD1S3IX count_2375__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i5.GSR = "ENABLED";
    FD1S3IX count_2375__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i6.GSR = "ENABLED";
    FD1S3IX count_2375__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i7.GSR = "ENABLED";
    FD1S3IX count_2375__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i8.GSR = "ENABLED";
    FD1S3IX count_2375__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i9.GSR = "ENABLED";
    FD1S3IX count_2375__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i10.GSR = "ENABLED";
    FD1S3IX count_2375__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i11.GSR = "ENABLED";
    FD1S3IX count_2375__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i12.GSR = "ENABLED";
    FD1S3IX count_2375__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i13.GSR = "ENABLED";
    FD1S3IX count_2375__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i14.GSR = "ENABLED";
    FD1S3IX count_2375__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i15.GSR = "ENABLED";
    FD1S3IX count_2375__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i16.GSR = "ENABLED";
    FD1S3IX count_2375__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i17.GSR = "ENABLED";
    FD1S3IX count_2375__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i18.GSR = "ENABLED";
    FD1S3IX count_2375__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i19.GSR = "ENABLED";
    FD1S3IX count_2375__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i20.GSR = "ENABLED";
    FD1S3IX count_2375__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i21.GSR = "ENABLED";
    FD1S3IX count_2375__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i22.GSR = "ENABLED";
    FD1S3IX count_2375__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i23.GSR = "ENABLED";
    FD1S3IX count_2375__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i24.GSR = "ENABLED";
    FD1S3IX count_2375__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i25.GSR = "ENABLED";
    FD1S3IX count_2375__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i26.GSR = "ENABLED";
    FD1S3IX count_2375__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i27.GSR = "ENABLED";
    FD1S3IX count_2375__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i28.GSR = "ENABLED";
    FD1S3IX count_2375__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i29.GSR = "ENABLED";
    FD1S3IX count_2375__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i30.GSR = "ENABLED";
    FD1S3IX count_2375__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28399), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2375__i31.GSR = "ENABLED";
    CCU2D sub_1883_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23817), .COUT(n23818));
    defparam sub_1883_add_2_11.INIT0 = 16'h5999;
    defparam sub_1883_add_2_11.INIT1 = 16'h5999;
    defparam sub_1883_add_2_11.INJECT1_0 = "NO";
    defparam sub_1883_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23816), .COUT(n23817));
    defparam sub_1883_add_2_9.INIT0 = 16'h5999;
    defparam sub_1883_add_2_9.INIT1 = 16'h5999;
    defparam sub_1883_add_2_9.INJECT1_0 = "NO";
    defparam sub_1883_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23819), .COUT(n23820));
    defparam sub_1883_add_2_15.INIT0 = 16'h5999;
    defparam sub_1883_add_2_15.INIT1 = 16'h5999;
    defparam sub_1883_add_2_15.INJECT1_0 = "NO";
    defparam sub_1883_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1881_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n23829));
    defparam sub_1881_add_2_1.INIT0 = 16'h0000;
    defparam sub_1881_add_2_1.INIT1 = 16'h5999;
    defparam sub_1881_add_2_1.INJECT1_0 = "NO";
    defparam sub_1881_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24100), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24099), .COUT(n24100), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24098), .COUT(n24099), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24097), .COUT(n24098), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24440), .S1(n7486));
    defparam sub_1884_add_2_33.INIT0 = 16'hf555;
    defparam sub_1884_add_2_33.INIT1 = 16'h0000;
    defparam sub_1884_add_2_33.INJECT1_0 = "NO";
    defparam sub_1884_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24096), .COUT(n24097), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24439), .COUT(n24440));
    defparam sub_1884_add_2_31.INIT0 = 16'hf555;
    defparam sub_1884_add_2_31.INIT1 = 16'hf555;
    defparam sub_1884_add_2_31.INJECT1_0 = "NO";
    defparam sub_1884_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24095), .COUT(n24096), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24438), .COUT(n24439));
    defparam sub_1884_add_2_29.INIT0 = 16'hf555;
    defparam sub_1884_add_2_29.INIT1 = 16'hf555;
    defparam sub_1884_add_2_29.INJECT1_0 = "NO";
    defparam sub_1884_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24437), .COUT(n24438));
    defparam sub_1884_add_2_27.INIT0 = 16'hf555;
    defparam sub_1884_add_2_27.INIT1 = 16'hf555;
    defparam sub_1884_add_2_27.INJECT1_0 = "NO";
    defparam sub_1884_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24436), .COUT(n24437));
    defparam sub_1884_add_2_25.INIT0 = 16'hf555;
    defparam sub_1884_add_2_25.INIT1 = 16'hf555;
    defparam sub_1884_add_2_25.INJECT1_0 = "NO";
    defparam sub_1884_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24094), .COUT(n24095), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24435), .COUT(n24436));
    defparam sub_1884_add_2_23.INIT0 = 16'hf555;
    defparam sub_1884_add_2_23.INIT1 = 16'hf555;
    defparam sub_1884_add_2_23.INJECT1_0 = "NO";
    defparam sub_1884_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24093), .COUT(n24094), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24092), .COUT(n24093), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24434), .COUT(n24435));
    defparam sub_1884_add_2_21.INIT0 = 16'hf555;
    defparam sub_1884_add_2_21.INIT1 = 16'hf555;
    defparam sub_1884_add_2_21.INJECT1_0 = "NO";
    defparam sub_1884_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24091), .COUT(n24092), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24090), .COUT(n24091), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24433), .COUT(n24434));
    defparam sub_1884_add_2_19.INIT0 = 16'hf555;
    defparam sub_1884_add_2_19.INIT1 = 16'hf555;
    defparam sub_1884_add_2_19.INJECT1_0 = "NO";
    defparam sub_1884_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24432), .COUT(n24433));
    defparam sub_1884_add_2_17.INIT0 = 16'hf555;
    defparam sub_1884_add_2_17.INIT1 = 16'hf555;
    defparam sub_1884_add_2_17.INJECT1_0 = "NO";
    defparam sub_1884_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24431), .COUT(n24432));
    defparam sub_1884_add_2_15.INIT0 = 16'hf555;
    defparam sub_1884_add_2_15.INIT1 = 16'hf555;
    defparam sub_1884_add_2_15.INJECT1_0 = "NO";
    defparam sub_1884_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24089), .COUT(n24090), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24088), .COUT(n24089), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24430), .COUT(n24431));
    defparam sub_1884_add_2_13.INIT0 = 16'hf555;
    defparam sub_1884_add_2_13.INIT1 = 16'hf555;
    defparam sub_1884_add_2_13.INJECT1_0 = "NO";
    defparam sub_1884_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24429), .COUT(n24430));
    defparam sub_1884_add_2_11.INIT0 = 16'hf555;
    defparam sub_1884_add_2_11.INIT1 = 16'hf555;
    defparam sub_1884_add_2_11.INJECT1_0 = "NO";
    defparam sub_1884_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24087), .COUT(n24088), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24428), .COUT(n24429));
    defparam sub_1884_add_2_9.INIT0 = 16'hf555;
    defparam sub_1884_add_2_9.INIT1 = 16'hf555;
    defparam sub_1884_add_2_9.INJECT1_0 = "NO";
    defparam sub_1884_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24427), .COUT(n24428));
    defparam sub_1884_add_2_7.INIT0 = 16'hf555;
    defparam sub_1884_add_2_7.INIT1 = 16'hf555;
    defparam sub_1884_add_2_7.INJECT1_0 = "NO";
    defparam sub_1884_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24426), .COUT(n24427));
    defparam sub_1884_add_2_5.INIT0 = 16'hf555;
    defparam sub_1884_add_2_5.INIT1 = 16'hf555;
    defparam sub_1884_add_2_5.INJECT1_0 = "NO";
    defparam sub_1884_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24086), .COUT(n24087), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24425), .COUT(n24426));
    defparam sub_1884_add_2_3.INIT0 = 16'hf555;
    defparam sub_1884_add_2_3.INIT1 = 16'hf555;
    defparam sub_1884_add_2_3.INJECT1_0 = "NO";
    defparam sub_1884_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1884_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24425));
    defparam sub_1884_add_2_1.INIT0 = 16'h0000;
    defparam sub_1884_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1884_add_2_1.INJECT1_0 = "NO";
    defparam sub_1884_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24085), .COUT(n24086), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24085), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23828), .S1(n7452));
    defparam sub_1883_add_2_33.INIT0 = 16'h5999;
    defparam sub_1883_add_2_33.INIT1 = 16'h0000;
    defparam sub_1883_add_2_33.INJECT1_0 = "NO";
    defparam sub_1883_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23827), .COUT(n23828));
    defparam sub_1883_add_2_31.INIT0 = 16'h5999;
    defparam sub_1883_add_2_31.INIT1 = 16'h5999;
    defparam sub_1883_add_2_31.INJECT1_0 = "NO";
    defparam sub_1883_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1883_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23826), .COUT(n23827));
    defparam sub_1883_add_2_29.INIT0 = 16'h5999;
    defparam sub_1883_add_2_29.INIT1 = 16'h5999;
    defparam sub_1883_add_2_29.INJECT1_0 = "NO";
    defparam sub_1883_add_2_29.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (GND_net, n7001, n28477, clk_255kHz, n6966, 
            n26942, n24743, n26945, n24741, debug_c_c, n241, n26947, 
            n24721, n2610, n26949, n24707, n26922, n12605, n26907, 
            n24716, n27027, n13534, n26939, n24755, n27025, n13535, 
            n27023, n13536, n27040, n13489, n27035, n13527) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n7001;
    input n28477;
    output clk_255kHz;
    output n6966;
    input n26942;
    output n24743;
    input n26945;
    output n24741;
    input debug_c_c;
    input n241;
    input n26947;
    output n24721;
    input n2610;
    input n26949;
    output n24707;
    input n26922;
    output n12605;
    input n26907;
    output n24716;
    input n27027;
    output n13534;
    input n26939;
    output n24755;
    input n27025;
    output n13535;
    input n27023;
    output n13536;
    input n27040;
    output n13489;
    input n27035;
    output n13527;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24408, n24407;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n24406, n24405, n24404, n24403, n24402, n24401, n24400, 
        n24399, n24398, n24397, n24396, n24395, n24394, n24393;
    wire [31:0]n134;
    
    wire n24491, n24490, n24489, n24488, n24487, n24486, n24485, 
        n24484, n24483, n24482, n24481, n24480, n24479, n24478, 
        n24477, n24264, n24263, n24262, n24261, n24260, n24259, 
        n24258, n24257, n24256, n24255, n24254, n24253, n24252, 
        n24251, n24250, n24249;
    
    CCU2D sub_1861_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24408), .S0(n7001));
    defparam sub_1861_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1861_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1861_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1861_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24407), .COUT(n24408));
    defparam sub_1861_add_2_32.INIT0 = 16'h5555;
    defparam sub_1861_add_2_32.INIT1 = 16'h5555;
    defparam sub_1861_add_2_32.INJECT1_0 = "NO";
    defparam sub_1861_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24406), .COUT(n24407));
    defparam sub_1861_add_2_30.INIT0 = 16'h5555;
    defparam sub_1861_add_2_30.INIT1 = 16'h5555;
    defparam sub_1861_add_2_30.INJECT1_0 = "NO";
    defparam sub_1861_add_2_30.INJECT1_1 = "NO";
    LUT4 i20344_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n26942), 
         .Z(n24743)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20344_2_lut_4_lut.init = 16'h1000;
    LUT4 i20347_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n26945), 
         .Z(n24741)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20347_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_1861_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24405), .COUT(n24406));
    defparam sub_1861_add_2_28.INIT0 = 16'h5555;
    defparam sub_1861_add_2_28.INIT1 = 16'h5555;
    defparam sub_1861_add_2_28.INJECT1_0 = "NO";
    defparam sub_1861_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24404), .COUT(n24405));
    defparam sub_1861_add_2_26.INIT0 = 16'h5555;
    defparam sub_1861_add_2_26.INIT1 = 16'h5555;
    defparam sub_1861_add_2_26.INJECT1_0 = "NO";
    defparam sub_1861_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24403), .COUT(n24404));
    defparam sub_1861_add_2_24.INIT0 = 16'h5555;
    defparam sub_1861_add_2_24.INIT1 = 16'h5555;
    defparam sub_1861_add_2_24.INJECT1_0 = "NO";
    defparam sub_1861_add_2_24.INJECT1_1 = "NO";
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=518, LSE_RLINE=521 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1861_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24402), .COUT(n24403));
    defparam sub_1861_add_2_22.INIT0 = 16'h5555;
    defparam sub_1861_add_2_22.INIT1 = 16'h5555;
    defparam sub_1861_add_2_22.INJECT1_0 = "NO";
    defparam sub_1861_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24401), .COUT(n24402));
    defparam sub_1861_add_2_20.INIT0 = 16'h5555;
    defparam sub_1861_add_2_20.INIT1 = 16'h5555;
    defparam sub_1861_add_2_20.INJECT1_0 = "NO";
    defparam sub_1861_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24400), .COUT(n24401));
    defparam sub_1861_add_2_18.INIT0 = 16'h5555;
    defparam sub_1861_add_2_18.INIT1 = 16'h5555;
    defparam sub_1861_add_2_18.INJECT1_0 = "NO";
    defparam sub_1861_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24399), .COUT(n24400));
    defparam sub_1861_add_2_16.INIT0 = 16'h5555;
    defparam sub_1861_add_2_16.INIT1 = 16'h5555;
    defparam sub_1861_add_2_16.INJECT1_0 = "NO";
    defparam sub_1861_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24398), .COUT(n24399));
    defparam sub_1861_add_2_14.INIT0 = 16'h5555;
    defparam sub_1861_add_2_14.INIT1 = 16'h5555;
    defparam sub_1861_add_2_14.INJECT1_0 = "NO";
    defparam sub_1861_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24397), .COUT(n24398));
    defparam sub_1861_add_2_12.INIT0 = 16'h5555;
    defparam sub_1861_add_2_12.INIT1 = 16'h5555;
    defparam sub_1861_add_2_12.INJECT1_0 = "NO";
    defparam sub_1861_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24396), .COUT(n24397));
    defparam sub_1861_add_2_10.INIT0 = 16'h5555;
    defparam sub_1861_add_2_10.INIT1 = 16'h5555;
    defparam sub_1861_add_2_10.INJECT1_0 = "NO";
    defparam sub_1861_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24395), .COUT(n24396));
    defparam sub_1861_add_2_8.INIT0 = 16'h5555;
    defparam sub_1861_add_2_8.INIT1 = 16'h5555;
    defparam sub_1861_add_2_8.INJECT1_0 = "NO";
    defparam sub_1861_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24394), .COUT(n24395));
    defparam sub_1861_add_2_6.INIT0 = 16'h5555;
    defparam sub_1861_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_1861_add_2_6.INJECT1_0 = "NO";
    defparam sub_1861_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24393), .COUT(n24394));
    defparam sub_1861_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1861_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_1861_add_2_4.INJECT1_0 = "NO";
    defparam sub_1861_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_1861_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24393));
    defparam sub_1861_add_2_2.INIT0 = 16'h0000;
    defparam sub_1861_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1861_add_2_2.INJECT1_0 = "NO";
    defparam sub_1861_add_2_2.INJECT1_1 = "NO";
    LUT4 i20349_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n26947), 
         .Z(n24721)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20349_2_lut_4_lut.init = 16'h1000;
    FD1S3IX count_2370__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2610), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i0.GSR = "ENABLED";
    LUT4 i20351_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n26949), 
         .Z(n24707)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20351_2_lut_4_lut.init = 16'h1000;
    LUT4 i20324_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n26922), 
         .Z(n12605)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20324_2_lut_4_lut.init = 16'h1000;
    LUT4 i20309_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n26907), 
         .Z(n24716)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20309_2_lut_4_lut.init = 16'h1000;
    LUT4 i20429_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n27027), 
         .Z(n13534)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20429_2_lut_4_lut.init = 16'h1000;
    LUT4 i20341_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n26939), 
         .Z(n24755)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20341_2_lut_4_lut.init = 16'h1000;
    LUT4 i20427_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n27025), 
         .Z(n13535)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20427_2_lut_4_lut.init = 16'h1000;
    LUT4 i20425_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n27023), 
         .Z(n13536)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20425_2_lut_4_lut.init = 16'h1000;
    LUT4 i20442_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n27040), 
         .Z(n13489)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20442_2_lut_4_lut.init = 16'h1000;
    CCU2D add_17800_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24491), 
          .S1(n6966));
    defparam add_17800_32.INIT0 = 16'h5555;
    defparam add_17800_32.INIT1 = 16'h0000;
    defparam add_17800_32.INJECT1_0 = "NO";
    defparam add_17800_32.INJECT1_1 = "NO";
    CCU2D add_17800_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24490), .COUT(n24491));
    defparam add_17800_30.INIT0 = 16'h5555;
    defparam add_17800_30.INIT1 = 16'h5555;
    defparam add_17800_30.INJECT1_0 = "NO";
    defparam add_17800_30.INJECT1_1 = "NO";
    CCU2D add_17800_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24489), .COUT(n24490));
    defparam add_17800_28.INIT0 = 16'h5555;
    defparam add_17800_28.INIT1 = 16'h5555;
    defparam add_17800_28.INJECT1_0 = "NO";
    defparam add_17800_28.INJECT1_1 = "NO";
    CCU2D add_17800_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24488), .COUT(n24489));
    defparam add_17800_26.INIT0 = 16'h5555;
    defparam add_17800_26.INIT1 = 16'h5555;
    defparam add_17800_26.INJECT1_0 = "NO";
    defparam add_17800_26.INJECT1_1 = "NO";
    CCU2D add_17800_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24487), .COUT(n24488));
    defparam add_17800_24.INIT0 = 16'h5555;
    defparam add_17800_24.INIT1 = 16'h5555;
    defparam add_17800_24.INJECT1_0 = "NO";
    defparam add_17800_24.INJECT1_1 = "NO";
    CCU2D add_17800_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24486), .COUT(n24487));
    defparam add_17800_22.INIT0 = 16'h5555;
    defparam add_17800_22.INIT1 = 16'h5555;
    defparam add_17800_22.INJECT1_0 = "NO";
    defparam add_17800_22.INJECT1_1 = "NO";
    CCU2D add_17800_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24485), .COUT(n24486));
    defparam add_17800_20.INIT0 = 16'h5555;
    defparam add_17800_20.INIT1 = 16'h5555;
    defparam add_17800_20.INJECT1_0 = "NO";
    defparam add_17800_20.INJECT1_1 = "NO";
    CCU2D add_17800_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24484), .COUT(n24485));
    defparam add_17800_18.INIT0 = 16'h5555;
    defparam add_17800_18.INIT1 = 16'h5555;
    defparam add_17800_18.INJECT1_0 = "NO";
    defparam add_17800_18.INJECT1_1 = "NO";
    CCU2D add_17800_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24483), .COUT(n24484));
    defparam add_17800_16.INIT0 = 16'h5555;
    defparam add_17800_16.INIT1 = 16'h5555;
    defparam add_17800_16.INJECT1_0 = "NO";
    defparam add_17800_16.INJECT1_1 = "NO";
    CCU2D add_17800_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24482), .COUT(n24483));
    defparam add_17800_14.INIT0 = 16'h5555;
    defparam add_17800_14.INIT1 = 16'h5555;
    defparam add_17800_14.INJECT1_0 = "NO";
    defparam add_17800_14.INJECT1_1 = "NO";
    CCU2D add_17800_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24481), .COUT(n24482));
    defparam add_17800_12.INIT0 = 16'h5555;
    defparam add_17800_12.INIT1 = 16'h5555;
    defparam add_17800_12.INJECT1_0 = "NO";
    defparam add_17800_12.INJECT1_1 = "NO";
    CCU2D add_17800_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24480), .COUT(n24481));
    defparam add_17800_10.INIT0 = 16'h5555;
    defparam add_17800_10.INIT1 = 16'h5555;
    defparam add_17800_10.INJECT1_0 = "NO";
    defparam add_17800_10.INJECT1_1 = "NO";
    CCU2D add_17800_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24479), 
          .COUT(n24480));
    defparam add_17800_8.INIT0 = 16'h5555;
    defparam add_17800_8.INIT1 = 16'h5555;
    defparam add_17800_8.INJECT1_0 = "NO";
    defparam add_17800_8.INJECT1_1 = "NO";
    CCU2D add_17800_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24478), 
          .COUT(n24479));
    defparam add_17800_6.INIT0 = 16'h5555;
    defparam add_17800_6.INIT1 = 16'h5555;
    defparam add_17800_6.INJECT1_0 = "NO";
    defparam add_17800_6.INJECT1_1 = "NO";
    CCU2D add_17800_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24477), 
          .COUT(n24478));
    defparam add_17800_4.INIT0 = 16'h5555;
    defparam add_17800_4.INIT1 = 16'h5aaa;
    defparam add_17800_4.INJECT1_0 = "NO";
    defparam add_17800_4.INJECT1_1 = "NO";
    FD1S3IX count_2370__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2610), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i1.GSR = "ENABLED";
    CCU2D add_17800_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24477));
    defparam add_17800_2.INIT0 = 16'h7000;
    defparam add_17800_2.INIT1 = 16'h5aaa;
    defparam add_17800_2.INJECT1_0 = "NO";
    defparam add_17800_2.INJECT1_1 = "NO";
    FD1S3IX count_2370__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2610), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i2.GSR = "ENABLED";
    FD1S3IX count_2370__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2610), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i3.GSR = "ENABLED";
    FD1S3IX count_2370__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2610), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i4.GSR = "ENABLED";
    FD1S3IX count_2370__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2610), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i5.GSR = "ENABLED";
    FD1S3IX count_2370__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2610), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i6.GSR = "ENABLED";
    FD1S3IX count_2370__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2610), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i7.GSR = "ENABLED";
    FD1S3IX count_2370__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2610), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i8.GSR = "ENABLED";
    FD1S3IX count_2370__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2610), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i9.GSR = "ENABLED";
    FD1S3IX count_2370__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i10.GSR = "ENABLED";
    FD1S3IX count_2370__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i11.GSR = "ENABLED";
    FD1S3IX count_2370__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i12.GSR = "ENABLED";
    FD1S3IX count_2370__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i13.GSR = "ENABLED";
    FD1S3IX count_2370__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i14.GSR = "ENABLED";
    FD1S3IX count_2370__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i15.GSR = "ENABLED";
    FD1S3IX count_2370__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i16.GSR = "ENABLED";
    FD1S3IX count_2370__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i17.GSR = "ENABLED";
    FD1S3IX count_2370__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i18.GSR = "ENABLED";
    FD1S3IX count_2370__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i19.GSR = "ENABLED";
    FD1S3IX count_2370__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i20.GSR = "ENABLED";
    FD1S3IX count_2370__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i21.GSR = "ENABLED";
    FD1S3IX count_2370__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i22.GSR = "ENABLED";
    FD1S3IX count_2370__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i23.GSR = "ENABLED";
    FD1S3IX count_2370__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i24.GSR = "ENABLED";
    FD1S3IX count_2370__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i25.GSR = "ENABLED";
    FD1S3IX count_2370__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i26.GSR = "ENABLED";
    FD1S3IX count_2370__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i27.GSR = "ENABLED";
    FD1S3IX count_2370__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i28.GSR = "ENABLED";
    FD1S3IX count_2370__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i29.GSR = "ENABLED";
    FD1S3IX count_2370__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i30.GSR = "ENABLED";
    FD1S3IX count_2370__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2610), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370__i31.GSR = "ENABLED";
    CCU2D count_2370_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24264), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_33.INIT1 = 16'h0000;
    defparam count_2370_add_4_33.INJECT1_0 = "NO";
    defparam count_2370_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24263), .COUT(n24264), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_31.INJECT1_0 = "NO";
    defparam count_2370_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24262), .COUT(n24263), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_29.INJECT1_0 = "NO";
    defparam count_2370_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24261), .COUT(n24262), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_27.INJECT1_0 = "NO";
    defparam count_2370_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24260), .COUT(n24261), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_25.INJECT1_0 = "NO";
    defparam count_2370_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24259), .COUT(n24260), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_23.INJECT1_0 = "NO";
    defparam count_2370_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24258), .COUT(n24259), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_21.INJECT1_0 = "NO";
    defparam count_2370_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24257), .COUT(n24258), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_19.INJECT1_0 = "NO";
    defparam count_2370_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24256), .COUT(n24257), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_17.INJECT1_0 = "NO";
    defparam count_2370_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24255), .COUT(n24256), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_15.INJECT1_0 = "NO";
    defparam count_2370_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24254), .COUT(n24255), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_13.INJECT1_0 = "NO";
    defparam count_2370_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24253), .COUT(n24254), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_11.INJECT1_0 = "NO";
    defparam count_2370_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24252), .COUT(n24253), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_9.INJECT1_0 = "NO";
    defparam count_2370_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24251), .COUT(n24252), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_7.INJECT1_0 = "NO";
    defparam count_2370_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24250), .COUT(n24251), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_5.INJECT1_0 = "NO";
    defparam count_2370_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24249), .COUT(n24250), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2370_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2370_add_4_3.INJECT1_0 = "NO";
    defparam count_2370_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2370_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24249), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2370_add_4_1.INIT0 = 16'hF000;
    defparam count_2370_add_4_1.INIT1 = 16'h0555;
    defparam count_2370_add_4_1.INJECT1_0 = "NO";
    defparam count_2370_add_4_1.INJECT1_1 = "NO";
    LUT4 i20437_2_lut_4_lut (.A(n28477), .B(clk_255kHz), .C(n6966), .D(n27035), 
         .Z(n13527)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i20437_2_lut_4_lut.init = 16'h1000;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (debug_c_c, n28414, n28477, databus, 
            n12647, n608, n610, \control_reg[7] , n12580, n10035, 
            Stepper_X_En_c, Stepper_X_Dir_c, n12583, Stepper_X_M2_c_2, 
            GND_net, Stepper_X_M1_c_1, \read_size[2] , n2615, n8336, 
            \steps_reg[7] , \register_addr[0] , \read_size[0] , n28425, 
            Stepper_X_M0_c_0, n579, limit_latched, prev_limit_latched, 
            prev_select, n28480, n3626, read_value, \register_addr[1] , 
            n19, limit_c_0, n12, VCC_net, Stepper_X_nFault_c, Stepper_X_Step_c, 
            n24815, n7140, n7174, n28401, n14714) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n28414;
    input n28477;
    input [31:0]databus;
    input n12647;
    input n608;
    input n610;
    output \control_reg[7] ;
    input n12580;
    input n10035;
    output Stepper_X_En_c;
    output Stepper_X_Dir_c;
    input n12583;
    output Stepper_X_M2_c_2;
    input GND_net;
    output Stepper_X_M1_c_1;
    output \read_size[2] ;
    input n2615;
    input n8336;
    output \steps_reg[7] ;
    input \register_addr[0] ;
    output \read_size[0] ;
    input n28425;
    output Stepper_X_M0_c_0;
    input n579;
    output limit_latched;
    output prev_limit_latched;
    output prev_select;
    input n28480;
    input n3626;
    output [31:0]read_value;
    input \register_addr[1] ;
    input n19;
    input limit_c_0;
    input n12;
    input VCC_net;
    input Stepper_X_nFault_c;
    output Stepper_X_Step_c;
    output n24815;
    output n7140;
    output n7174;
    input n28401;
    input n14714;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n24212;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n224;
    
    wire n24211, n24210, n24209, n24208;
    wire [31:0]n3627;
    
    wire n1, n2, n24207, n24206, n24205, prev_step_clk, step_clk, 
        n182, n24204, n1_adj_1, n2_adj_2, n26828, n26826, n26827, 
        n1_adj_3, n2_adj_4, n24203;
    wire [31:0]n100;
    
    wire n26864, n26834, n24202, n1_adj_5, n24201, n24200, n24199, 
        n24198, n16939;
    wire [31:0]n99;
    
    wire n24197, n26832, n26833, n26862, n26863, n28412, fault_latched, 
        n11, n17997, int_step, n49, n62_adj_6, n58_adj_7, n50_adj_8, 
        n41, n60, n54_adj_9, n42_adj_10, n52_adj_11, n38_adj_12, 
        n56_adj_13, n46_adj_14;
    
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n28414), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n28414), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n28414), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n28414), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n28414), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n28414), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n28414), .PD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n12647), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12647), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n12580), .CD(n10035), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n12580), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n12580), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n12583), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n12580), .PD(n28477), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n12583), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24212), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n12580), .PD(n28477), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n8336), .SP(n2615), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24211), .COUT(n24212), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24210), .COUT(n24211), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24209), .COUT(n24210), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24208), .COUT(n24209), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    FD1S3IX steps_reg__i31 (.D(n3627[31]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3627[30]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3627[29]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3627[28]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3627[27]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3627[26]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3627[25]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3627[24]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3627[23]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3627[22]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3627[21]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3627[20]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3627[19]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3627[18]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3627[17]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3627[16]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3627[15]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3627[14]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3627[13]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3627[12]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3627[11]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3627[10]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3627[9]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3627[8]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3627[7]), .CK(debug_c_c), .CD(n28477), 
            .Q(\steps_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3627[6]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3627[5]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3627[4]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3627[3]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3627[2]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3627[1]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i13400_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13400_2_lut.init = 16'h2222;
    LUT4 i10937_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i10937_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24207), .COUT(n24208), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24206), .COUT(n24207), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    FD1S3IX steps_reg__i0 (.D(n3627[0]), .CK(debug_c_c), .CD(n28477), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n28425), .SP(n2615), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24205), .COUT(n24206), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12583), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12647), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n28480), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24204), .COUT(n24205), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    LUT4 i13399_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13399_2_lut.init = 16'h2222;
    LUT4 mux_1735_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2_adj_2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1735_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3626), 
         .Z(n3627[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i32_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n26828), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    PFUMX i20132 (.BLUT(n26826), .ALUT(n26827), .C0(\register_addr[1] ), 
          .Z(n26828));
    LUT4 i13398_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_3)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13398_2_lut.init = 16'h2222;
    LUT4 mux_1517_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3626), .Z(n3627[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i1_3_lut.init = 16'hcaca;
    LUT4 i10938_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n2_adj_4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i10938_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24203), .COUT(n24204), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n26864), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n26834), .SP(n2615), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24202), .COUT(n24203), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    LUT4 i13397_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_5)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13397_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24201), .COUT(n24202), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(\steps_reg[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24200), .COUT(n24201), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24199), .COUT(n24200), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24198), .COUT(n24199), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 i10940_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n16939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i10940_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[18]), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n99[18])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'ha088;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24197), .COUT(n24198), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n19), .D1(prev_step_clk), 
          .COUT(n24197), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_1517_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3626), 
         .Z(n3627[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i22_3_lut.init = 16'hcaca;
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    PFUMX i20138 (.BLUT(n26832), .ALUT(n26833), .C0(\register_addr[1] ), 
          .Z(n26834));
    LUT4 mux_1517_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3626), 
         .Z(n3627[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3626), 
         .Z(n3627[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i11_3_lut.init = 16'hcaca;
    PFUMX mux_1735_Mux_3_i3 (.BLUT(n1), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    LUT4 mux_1517_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3626), .Z(n3627[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i10_3_lut.init = 16'hcaca;
    PFUMX mux_1735_Mux_4_i3 (.BLUT(n1_adj_1), .ALUT(n2_adj_2), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1735_Mux_5_i3 (.BLUT(n1_adj_3), .ALUT(n2_adj_4), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    LUT4 mux_1517_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3626), .Z(n3627[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3626), .Z(n3627[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3626), .Z(n3627[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3626), .Z(n3627[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3626), .Z(n3627[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i5_3_lut.init = 16'hcaca;
    PFUMX mux_1735_Mux_6_i3 (.BLUT(n1_adj_5), .ALUT(n16939), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    FD1P3AX read_value__i18 (.D(n99[18]), .SP(n2615), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    LUT4 mux_1517_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3626), .Z(n3627[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3626), .Z(n3627[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3626), .Z(n3627[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i2_3_lut.init = 16'hcaca;
    PFUMX i20168 (.BLUT(n26862), .ALUT(n26863), .C0(\register_addr[0] ), 
          .Z(n26864));
    LUT4 i2_3_lut_rep_291 (.A(prev_step_clk), .B(n19), .C(step_clk), .Z(n28412)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i2_3_lut_rep_291.init = 16'h4040;
    LUT4 i20136_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n26832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20136_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3626), 
         .Z(n3627[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i31_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut (.A(prev_step_clk), .B(n19), .C(step_clk), .D(n28477), 
         .Z(n11)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_4_lut.init = 16'h004a;
    LUT4 i20166_3_lut (.A(Stepper_X_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n26862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20166_3_lut.init = 16'hcaca;
    LUT4 i20167_3_lut (.A(n19), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n26863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20167_3_lut.init = 16'hcaca;
    LUT4 i20130_3_lut (.A(Stepper_X_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n26826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20130_3_lut.init = 16'hcaca;
    LUT4 i20131_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n26827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20131_3_lut.init = 16'hcaca;
    LUT4 i20137_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n26833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20137_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3626), 
         .Z(n3627[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3626), 
         .Z(n3627[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i21_3_lut.init = 16'hcaca;
    LUT4 i13618_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13618_4_lut.init = 16'hc088;
    LUT4 i13619_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13619_4_lut.init = 16'hc088;
    LUT4 i13620_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13620_4_lut.init = 16'hc088;
    LUT4 i13621_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13621_4_lut.init = 16'hc088;
    LUT4 i13622_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13622_4_lut.init = 16'hc088;
    LUT4 i13623_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13623_4_lut.init = 16'hc088;
    PFUMX i12011 (.BLUT(n17997), .ALUT(n12), .C0(\register_addr[0] ), 
          .Z(n100[7]));
    LUT4 mux_1517_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3626), 
         .Z(n3627[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i29_3_lut.init = 16'hcaca;
    LUT4 i13624_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13624_4_lut.init = 16'hc088;
    LUT4 i13625_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13625_4_lut.init = 16'hc088;
    LUT4 i13626_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13626_4_lut.init = 16'hc088;
    LUT4 i13627_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13627_4_lut.init = 16'hc088;
    LUT4 i13628_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13628_4_lut.init = 16'hc088;
    LUT4 i13629_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13629_4_lut.init = 16'hc088;
    LUT4 i13630_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13630_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_1 (.A(\register_addr[1] ), .B(div_factor_reg[17]), 
         .C(steps_reg[17]), .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_1.init = 16'ha088;
    LUT4 i13631_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13631_4_lut.init = 16'hc088;
    LUT4 i13632_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13632_4_lut.init = 16'hc088;
    LUT4 i13633_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13633_4_lut.init = 16'hc088;
    LUT4 i13634_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13634_4_lut.init = 16'hc088;
    LUT4 i13635_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13635_4_lut.init = 16'hc088;
    LUT4 i13636_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13636_4_lut.init = 16'hc088;
    LUT4 i13637_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13637_4_lut.init = 16'hc088;
    LUT4 i13638_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13638_4_lut.init = 16'hc088;
    LUT4 i13639_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13639_4_lut.init = 16'hc088;
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    LUT4 mux_1517_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3626), 
         .Z(n3627[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i28_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1517_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3626), 
         .Z(n3627[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3626), 
         .Z(n3627[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i20_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n28412), .SP(n11), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12647), .CD(n28477), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    LUT4 mux_1517_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3626), 
         .Z(n3627[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3626), 
         .Z(n3627[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3626), 
         .Z(n3627[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i14_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_6), .C(n58_adj_7), .D(n50_adj_8), 
         .Z(n24815)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 mux_1517_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3626), 
         .Z(n3627[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3626), 
         .Z(n3627[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i13_3_lut.init = 16'hcaca;
    LUT4 i17_4_lut (.A(steps_reg[12]), .B(steps_reg[18]), .C(steps_reg[17]), 
         .D(steps_reg[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54_adj_9), .D(n42_adj_10), 
         .Z(n62_adj_6)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[28]), .B(n52_adj_11), .C(n38_adj_12), 
         .D(steps_reg[24]), .Z(n58_adj_7)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[11]), .B(steps_reg[6]), .C(steps_reg[3]), 
         .D(steps_reg[9]), .Z(n50_adj_8)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[26]), .B(steps_reg[0]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[22]), .B(n56_adj_13), .C(n46_adj_14), 
         .D(steps_reg[1]), .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 mux_1517_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3626), 
         .Z(n3627[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3626), 
         .Z(n3627[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3626), 
         .Z(n3627[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i17_3_lut.init = 16'hcaca;
    LUT4 i22_4_lut (.A(steps_reg[15]), .B(steps_reg[14]), .C(steps_reg[23]), 
         .D(steps_reg[19]), .Z(n54_adj_9)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 mux_1517_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3626), 
         .Z(n3627[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i24_3_lut.init = 16'hcaca;
    LUT4 i10_2_lut (.A(steps_reg[20]), .B(steps_reg[29]), .Z(n42_adj_10)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[31]), .B(steps_reg[2]), .C(steps_reg[13]), 
         .D(steps_reg[4]), .Z(n56_adj_13)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 mux_1517_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3626), 
         .Z(n3627[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i16_3_lut.init = 16'hcaca;
    LUT4 i14_2_lut (.A(steps_reg[8]), .B(steps_reg[16]), .Z(n46_adj_14)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[5]), .B(steps_reg[21]), .C(steps_reg[27]), 
         .D(steps_reg[25]), .Z(n52_adj_11)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i12009_3_lut (.A(\control_reg[7] ), .B(div_factor_reg[7]), .C(\register_addr[1] ), 
         .Z(n17997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i12009_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut (.A(steps_reg[30]), .B(\steps_reg[7] ), .Z(n38_adj_12)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1517_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3626), 
         .Z(n3627[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1517_i23_3_lut.init = 16'hcaca;
    ClockDivider_U7 step_clk_gen (.GND_net(GND_net), .n7140(n7140), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n28477(n28477), .div_factor_reg({div_factor_reg}), 
            .n7174(n7174), .n28401(n28401), .n14714(n14714)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (GND_net, n7140, step_clk, debug_c_c, n28477, 
            div_factor_reg, n7174, n28401, n14714) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n7140;
    output step_clk;
    input debug_c_c;
    input n28477;
    input [31:0]div_factor_reg;
    output n7174;
    input n28401;
    input n14714;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n23992;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n23993, n23991, n23990, n23989, n23988;
    wire [31:0]n40;
    
    wire n23987, n23986, n23985, n23984, n23983, n23982, n23981, 
        n23980, n23979, n23978, n23977, n7105, n23976, n23975, 
        n23974, n23973, n23972;
    wire [31:0]n134;
    
    wire n23971, n23970, n23969, n23968, n23967, n23966, n23965, 
        n23964, n23963, n24328, n24327, n24326, n23962, n24325, 
        n24324, n24323, n24322, n24321, n23961, n24320, n24319, 
        n24318, n24317, n24316, n24315, n24314, n24313, n23960, 
        n23959, n23958, n23957, n24148, n24147, n24146, n24145, 
        n24144, n24143, n24142, n24141, n24140, n24139, n24138, 
        n24137, n24136, n24135, n24134, n24133, n24004, n24003, 
        n24002, n24001, n24000, n23999, n23998, n23997, n23996, 
        n23995, n23994;
    
    CCU2D sub_1866_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23992), .COUT(n23993));
    defparam sub_1866_add_2_9.INIT0 = 16'h5999;
    defparam sub_1866_add_2_9.INIT1 = 16'h5999;
    defparam sub_1866_add_2_9.INJECT1_0 = "NO";
    defparam sub_1866_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23991), .COUT(n23992));
    defparam sub_1866_add_2_7.INIT0 = 16'h5999;
    defparam sub_1866_add_2_7.INIT1 = 16'h5999;
    defparam sub_1866_add_2_7.INJECT1_0 = "NO";
    defparam sub_1866_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23990), .COUT(n23991));
    defparam sub_1866_add_2_5.INIT0 = 16'h5999;
    defparam sub_1866_add_2_5.INIT1 = 16'h5999;
    defparam sub_1866_add_2_5.INJECT1_0 = "NO";
    defparam sub_1866_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23989), .COUT(n23990));
    defparam sub_1866_add_2_3.INIT0 = 16'h5999;
    defparam sub_1866_add_2_3.INIT1 = 16'h5999;
    defparam sub_1866_add_2_3.INJECT1_0 = "NO";
    defparam sub_1866_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n23989));
    defparam sub_1866_add_2_1.INIT0 = 16'h0000;
    defparam sub_1866_add_2_1.INIT1 = 16'h5999;
    defparam sub_1866_add_2_1.INJECT1_0 = "NO";
    defparam sub_1866_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23988), .S1(n7140));
    defparam sub_1868_add_2_33.INIT0 = 16'h5999;
    defparam sub_1868_add_2_33.INIT1 = 16'h0000;
    defparam sub_1868_add_2_33.INJECT1_0 = "NO";
    defparam sub_1868_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23987), .COUT(n23988));
    defparam sub_1868_add_2_31.INIT0 = 16'h5999;
    defparam sub_1868_add_2_31.INIT1 = 16'h5999;
    defparam sub_1868_add_2_31.INJECT1_0 = "NO";
    defparam sub_1868_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23986), .COUT(n23987));
    defparam sub_1868_add_2_29.INIT0 = 16'h5999;
    defparam sub_1868_add_2_29.INIT1 = 16'h5999;
    defparam sub_1868_add_2_29.INJECT1_0 = "NO";
    defparam sub_1868_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23985), .COUT(n23986));
    defparam sub_1868_add_2_27.INIT0 = 16'h5999;
    defparam sub_1868_add_2_27.INIT1 = 16'h5999;
    defparam sub_1868_add_2_27.INJECT1_0 = "NO";
    defparam sub_1868_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23984), .COUT(n23985));
    defparam sub_1868_add_2_25.INIT0 = 16'h5999;
    defparam sub_1868_add_2_25.INIT1 = 16'h5999;
    defparam sub_1868_add_2_25.INJECT1_0 = "NO";
    defparam sub_1868_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23983), .COUT(n23984));
    defparam sub_1868_add_2_23.INIT0 = 16'h5999;
    defparam sub_1868_add_2_23.INIT1 = 16'h5999;
    defparam sub_1868_add_2_23.INJECT1_0 = "NO";
    defparam sub_1868_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23982), .COUT(n23983));
    defparam sub_1868_add_2_21.INIT0 = 16'h5999;
    defparam sub_1868_add_2_21.INIT1 = 16'h5999;
    defparam sub_1868_add_2_21.INJECT1_0 = "NO";
    defparam sub_1868_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23981), .COUT(n23982));
    defparam sub_1868_add_2_19.INIT0 = 16'h5999;
    defparam sub_1868_add_2_19.INIT1 = 16'h5999;
    defparam sub_1868_add_2_19.INJECT1_0 = "NO";
    defparam sub_1868_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23980), .COUT(n23981));
    defparam sub_1868_add_2_17.INIT0 = 16'h5999;
    defparam sub_1868_add_2_17.INIT1 = 16'h5999;
    defparam sub_1868_add_2_17.INJECT1_0 = "NO";
    defparam sub_1868_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23979), .COUT(n23980));
    defparam sub_1868_add_2_15.INIT0 = 16'h5999;
    defparam sub_1868_add_2_15.INIT1 = 16'h5999;
    defparam sub_1868_add_2_15.INJECT1_0 = "NO";
    defparam sub_1868_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23978), .COUT(n23979));
    defparam sub_1868_add_2_13.INIT0 = 16'h5999;
    defparam sub_1868_add_2_13.INIT1 = 16'h5999;
    defparam sub_1868_add_2_13.INJECT1_0 = "NO";
    defparam sub_1868_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23977), .COUT(n23978));
    defparam sub_1868_add_2_11.INIT0 = 16'h5999;
    defparam sub_1868_add_2_11.INIT1 = 16'h5999;
    defparam sub_1868_add_2_11.INJECT1_0 = "NO";
    defparam sub_1868_add_2_11.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7105), .CK(debug_c_c), .CD(n28477), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1868_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23976), .COUT(n23977));
    defparam sub_1868_add_2_9.INIT0 = 16'h5999;
    defparam sub_1868_add_2_9.INIT1 = 16'h5999;
    defparam sub_1868_add_2_9.INJECT1_0 = "NO";
    defparam sub_1868_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23975), .COUT(n23976));
    defparam sub_1868_add_2_7.INIT0 = 16'h5999;
    defparam sub_1868_add_2_7.INIT1 = 16'h5999;
    defparam sub_1868_add_2_7.INJECT1_0 = "NO";
    defparam sub_1868_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23974), .COUT(n23975));
    defparam sub_1868_add_2_5.INIT0 = 16'h5999;
    defparam sub_1868_add_2_5.INIT1 = 16'h5999;
    defparam sub_1868_add_2_5.INJECT1_0 = "NO";
    defparam sub_1868_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n23973), .COUT(n23974));
    defparam sub_1868_add_2_3.INIT0 = 16'h5999;
    defparam sub_1868_add_2_3.INIT1 = 16'h5999;
    defparam sub_1868_add_2_3.INJECT1_0 = "NO";
    defparam sub_1868_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1868_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n23973));
    defparam sub_1868_add_2_1.INIT0 = 16'h0000;
    defparam sub_1868_add_2_1.INIT1 = 16'h5999;
    defparam sub_1868_add_2_1.INJECT1_0 = "NO";
    defparam sub_1868_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23972), .S1(n7174));
    defparam sub_1869_add_2_33.INIT0 = 16'hf555;
    defparam sub_1869_add_2_33.INIT1 = 16'h0000;
    defparam sub_1869_add_2_33.INJECT1_0 = "NO";
    defparam sub_1869_add_2_33.INJECT1_1 = "NO";
    FD1S3IX count_2372__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i0.GSR = "ENABLED";
    CCU2D sub_1869_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23971), .COUT(n23972));
    defparam sub_1869_add_2_31.INIT0 = 16'hf555;
    defparam sub_1869_add_2_31.INIT1 = 16'hf555;
    defparam sub_1869_add_2_31.INJECT1_0 = "NO";
    defparam sub_1869_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23970), .COUT(n23971));
    defparam sub_1869_add_2_29.INIT0 = 16'hf555;
    defparam sub_1869_add_2_29.INIT1 = 16'hf555;
    defparam sub_1869_add_2_29.INJECT1_0 = "NO";
    defparam sub_1869_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23969), .COUT(n23970));
    defparam sub_1869_add_2_27.INIT0 = 16'hf555;
    defparam sub_1869_add_2_27.INIT1 = 16'hf555;
    defparam sub_1869_add_2_27.INJECT1_0 = "NO";
    defparam sub_1869_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23968), .COUT(n23969));
    defparam sub_1869_add_2_25.INIT0 = 16'hf555;
    defparam sub_1869_add_2_25.INIT1 = 16'hf555;
    defparam sub_1869_add_2_25.INJECT1_0 = "NO";
    defparam sub_1869_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23967), .COUT(n23968));
    defparam sub_1869_add_2_23.INIT0 = 16'hf555;
    defparam sub_1869_add_2_23.INIT1 = 16'hf555;
    defparam sub_1869_add_2_23.INJECT1_0 = "NO";
    defparam sub_1869_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23966), .COUT(n23967));
    defparam sub_1869_add_2_21.INIT0 = 16'hf555;
    defparam sub_1869_add_2_21.INIT1 = 16'hf555;
    defparam sub_1869_add_2_21.INJECT1_0 = "NO";
    defparam sub_1869_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23965), .COUT(n23966));
    defparam sub_1869_add_2_19.INIT0 = 16'hf555;
    defparam sub_1869_add_2_19.INIT1 = 16'hf555;
    defparam sub_1869_add_2_19.INJECT1_0 = "NO";
    defparam sub_1869_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23964), .COUT(n23965));
    defparam sub_1869_add_2_17.INIT0 = 16'hf555;
    defparam sub_1869_add_2_17.INIT1 = 16'hf555;
    defparam sub_1869_add_2_17.INJECT1_0 = "NO";
    defparam sub_1869_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23963), .COUT(n23964));
    defparam sub_1869_add_2_15.INIT0 = 16'hf555;
    defparam sub_1869_add_2_15.INIT1 = 16'hf555;
    defparam sub_1869_add_2_15.INJECT1_0 = "NO";
    defparam sub_1869_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24328), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_33.INIT1 = 16'h0000;
    defparam count_2372_add_4_33.INJECT1_0 = "NO";
    defparam count_2372_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24327), .COUT(n24328), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_31.INJECT1_0 = "NO";
    defparam count_2372_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24326), .COUT(n24327), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_29.INJECT1_0 = "NO";
    defparam count_2372_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23962), .COUT(n23963));
    defparam sub_1869_add_2_13.INIT0 = 16'hf555;
    defparam sub_1869_add_2_13.INIT1 = 16'hf555;
    defparam sub_1869_add_2_13.INJECT1_0 = "NO";
    defparam sub_1869_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24325), .COUT(n24326), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_27.INJECT1_0 = "NO";
    defparam count_2372_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24324), .COUT(n24325), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_25.INJECT1_0 = "NO";
    defparam count_2372_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24323), .COUT(n24324), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_23.INJECT1_0 = "NO";
    defparam count_2372_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24322), .COUT(n24323), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_21.INJECT1_0 = "NO";
    defparam count_2372_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24321), .COUT(n24322), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_19.INJECT1_0 = "NO";
    defparam count_2372_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23961), .COUT(n23962));
    defparam sub_1869_add_2_11.INIT0 = 16'hf555;
    defparam sub_1869_add_2_11.INIT1 = 16'hf555;
    defparam sub_1869_add_2_11.INJECT1_0 = "NO";
    defparam sub_1869_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24320), .COUT(n24321), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_17.INJECT1_0 = "NO";
    defparam count_2372_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24319), .COUT(n24320), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_15.INJECT1_0 = "NO";
    defparam count_2372_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24318), .COUT(n24319), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_13.INJECT1_0 = "NO";
    defparam count_2372_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24317), .COUT(n24318), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_11.INJECT1_0 = "NO";
    defparam count_2372_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24316), .COUT(n24317), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_9.INJECT1_0 = "NO";
    defparam count_2372_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24315), .COUT(n24316), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_7.INJECT1_0 = "NO";
    defparam count_2372_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24314), .COUT(n24315), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_5.INJECT1_0 = "NO";
    defparam count_2372_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24313), .COUT(n24314), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2372_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2372_add_4_3.INJECT1_0 = "NO";
    defparam count_2372_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2372_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24313), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372_add_4_1.INIT0 = 16'hF000;
    defparam count_2372_add_4_1.INIT1 = 16'h0555;
    defparam count_2372_add_4_1.INJECT1_0 = "NO";
    defparam count_2372_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23960), .COUT(n23961));
    defparam sub_1869_add_2_9.INIT0 = 16'hf555;
    defparam sub_1869_add_2_9.INIT1 = 16'hf555;
    defparam sub_1869_add_2_9.INJECT1_0 = "NO";
    defparam sub_1869_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23959), .COUT(n23960));
    defparam sub_1869_add_2_7.INIT0 = 16'hf555;
    defparam sub_1869_add_2_7.INIT1 = 16'hf555;
    defparam sub_1869_add_2_7.INJECT1_0 = "NO";
    defparam sub_1869_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23958), .COUT(n23959));
    defparam sub_1869_add_2_5.INIT0 = 16'hf555;
    defparam sub_1869_add_2_5.INIT1 = 16'hf555;
    defparam sub_1869_add_2_5.INJECT1_0 = "NO";
    defparam sub_1869_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23957), .COUT(n23958));
    defparam sub_1869_add_2_3.INIT0 = 16'hf555;
    defparam sub_1869_add_2_3.INIT1 = 16'hf555;
    defparam sub_1869_add_2_3.INJECT1_0 = "NO";
    defparam sub_1869_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24148), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24147), .COUT(n24148), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1869_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n23957));
    defparam sub_1869_add_2_1.INIT0 = 16'h0000;
    defparam sub_1869_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1869_add_2_1.INJECT1_0 = "NO";
    defparam sub_1869_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24146), .COUT(n24147), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24145), .COUT(n24146), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24144), .COUT(n24145), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24143), .COUT(n24144), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24142), .COUT(n24143), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24141), .COUT(n24142), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24140), .COUT(n24141), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24139), .COUT(n24140), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24138), .COUT(n24139), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24137), .COUT(n24138), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24136), .COUT(n24137), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24135), .COUT(n24136), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24134), .COUT(n24135), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24133), .COUT(n24134), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24133), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28401), .PD(n14714), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28401), .CD(n14714), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1S3IX count_2372__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i1.GSR = "ENABLED";
    FD1S3IX count_2372__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i2.GSR = "ENABLED";
    FD1S3IX count_2372__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i3.GSR = "ENABLED";
    FD1S3IX count_2372__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i4.GSR = "ENABLED";
    FD1S3IX count_2372__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i5.GSR = "ENABLED";
    FD1S3IX count_2372__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i6.GSR = "ENABLED";
    FD1S3IX count_2372__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i7.GSR = "ENABLED";
    FD1S3IX count_2372__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i8.GSR = "ENABLED";
    FD1S3IX count_2372__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i9.GSR = "ENABLED";
    FD1S3IX count_2372__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i10.GSR = "ENABLED";
    FD1S3IX count_2372__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i11.GSR = "ENABLED";
    FD1S3IX count_2372__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i12.GSR = "ENABLED";
    FD1S3IX count_2372__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i13.GSR = "ENABLED";
    FD1S3IX count_2372__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i14.GSR = "ENABLED";
    FD1S3IX count_2372__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i15.GSR = "ENABLED";
    FD1S3IX count_2372__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i16.GSR = "ENABLED";
    FD1S3IX count_2372__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i17.GSR = "ENABLED";
    FD1S3IX count_2372__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i18.GSR = "ENABLED";
    FD1S3IX count_2372__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i19.GSR = "ENABLED";
    FD1S3IX count_2372__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i20.GSR = "ENABLED";
    FD1S3IX count_2372__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i21.GSR = "ENABLED";
    FD1S3IX count_2372__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i22.GSR = "ENABLED";
    FD1S3IX count_2372__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i23.GSR = "ENABLED";
    FD1S3IX count_2372__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i24.GSR = "ENABLED";
    FD1S3IX count_2372__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i25.GSR = "ENABLED";
    FD1S3IX count_2372__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i26.GSR = "ENABLED";
    FD1S3IX count_2372__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i27.GSR = "ENABLED";
    FD1S3IX count_2372__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i28.GSR = "ENABLED";
    FD1S3IX count_2372__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i29.GSR = "ENABLED";
    FD1S3IX count_2372__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i30.GSR = "ENABLED";
    FD1S3IX count_2372__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28401), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2372__i31.GSR = "ENABLED";
    CCU2D sub_1866_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24004), .S1(n7105));
    defparam sub_1866_add_2_33.INIT0 = 16'h5555;
    defparam sub_1866_add_2_33.INIT1 = 16'h0000;
    defparam sub_1866_add_2_33.INJECT1_0 = "NO";
    defparam sub_1866_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24003), .COUT(n24004));
    defparam sub_1866_add_2_31.INIT0 = 16'h5999;
    defparam sub_1866_add_2_31.INIT1 = 16'h5999;
    defparam sub_1866_add_2_31.INJECT1_0 = "NO";
    defparam sub_1866_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24002), .COUT(n24003));
    defparam sub_1866_add_2_29.INIT0 = 16'h5999;
    defparam sub_1866_add_2_29.INIT1 = 16'h5999;
    defparam sub_1866_add_2_29.INJECT1_0 = "NO";
    defparam sub_1866_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24001), .COUT(n24002));
    defparam sub_1866_add_2_27.INIT0 = 16'h5999;
    defparam sub_1866_add_2_27.INIT1 = 16'h5999;
    defparam sub_1866_add_2_27.INJECT1_0 = "NO";
    defparam sub_1866_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24000), .COUT(n24001));
    defparam sub_1866_add_2_25.INIT0 = 16'h5999;
    defparam sub_1866_add_2_25.INIT1 = 16'h5999;
    defparam sub_1866_add_2_25.INJECT1_0 = "NO";
    defparam sub_1866_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23999), .COUT(n24000));
    defparam sub_1866_add_2_23.INIT0 = 16'h5999;
    defparam sub_1866_add_2_23.INIT1 = 16'h5999;
    defparam sub_1866_add_2_23.INJECT1_0 = "NO";
    defparam sub_1866_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23998), .COUT(n23999));
    defparam sub_1866_add_2_21.INIT0 = 16'h5999;
    defparam sub_1866_add_2_21.INIT1 = 16'h5999;
    defparam sub_1866_add_2_21.INJECT1_0 = "NO";
    defparam sub_1866_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23997), .COUT(n23998));
    defparam sub_1866_add_2_19.INIT0 = 16'h5999;
    defparam sub_1866_add_2_19.INIT1 = 16'h5999;
    defparam sub_1866_add_2_19.INJECT1_0 = "NO";
    defparam sub_1866_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23996), .COUT(n23997));
    defparam sub_1866_add_2_17.INIT0 = 16'h5999;
    defparam sub_1866_add_2_17.INIT1 = 16'h5999;
    defparam sub_1866_add_2_17.INJECT1_0 = "NO";
    defparam sub_1866_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23995), .COUT(n23996));
    defparam sub_1866_add_2_15.INIT0 = 16'h5999;
    defparam sub_1866_add_2_15.INIT1 = 16'h5999;
    defparam sub_1866_add_2_15.INJECT1_0 = "NO";
    defparam sub_1866_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23994), .COUT(n23995));
    defparam sub_1866_add_2_13.INIT0 = 16'h5999;
    defparam sub_1866_add_2_13.INIT1 = 16'h5999;
    defparam sub_1866_add_2_13.INJECT1_0 = "NO";
    defparam sub_1866_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1866_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23993), .COUT(n23994));
    defparam sub_1866_add_2_11.INIT0 = 16'h5999;
    defparam sub_1866_add_2_11.INIT1 = 16'h5999;
    defparam sub_1866_add_2_11.INJECT1_0 = "NO";
    defparam sub_1866_add_2_11.INJECT1_1 = "NO";
    
endmodule
