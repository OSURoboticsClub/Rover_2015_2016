// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Mon Jan 18 19:32:23 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    output expansion4 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    
    wire GND_net, VCC_net, n9396_c, n9395, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, signal_light_c, rc_ch1_c, rc_ch2_c, rc_ch3_c, rc_ch4_c, 
        rc_ch7_c, rc_ch8_c, xbee_pause_c, debug_c_7, debug_c_5, debug_c_4, 
        debug_c_3, debug_c_2;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire rw, n28352;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    
    wire n14473, n32404, n32403, n28360, n20528, n12620, n12434, 
        n14446, n31582, n10513, n1;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n31033, n27793, n27792, n4, n31025, n2, n27791, n27790, 
        n32400, n6, n28386, n27789;
    wire [31:0]n1286;
    
    wire n27788, n27787, n28331, n6_adj_393, n183, n2_adj_394, n11753;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[12:21])
    
    wire n12224;
    wire [7:0]n7893;
    
    wire n9, n11645, n1_adj_395, n32396, n32395, n15, n2_adj_396, 
        n30934, n18, n9633, n30, n241;
    wire [7:0]read_value_adj_688;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(63[12:22])
    wire [2:0]read_size_adj_689;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(64[12:21])
    
    wire n64;
    wire [15:0]n281;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]read_value_adj_693;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_694;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select, n6_adj_439, n15_adj_440, n3363;
    wire [31:0]n224;
    
    wire n2_adj_442, n302;
    wire [31:0]n3451;
    wire [7:0]n571;
    
    wire n14322;
    wire [31:0]n580;
    
    wire n12138;
    wire [7:0]control_reg_adj_702;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_704;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping;
    wire [31:0]read_value_adj_705;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_706;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_478, n52, n4_adj_479, n7912, n19896;
    wire [7:0]control_reg_adj_742;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_744;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping_adj_483;
    wire [31:0]read_value_adj_745;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_746;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_518, n30999, n30363;
    wire [31:0]n3181;
    
    wire n3589, n12098, n30283, n16, motor_pwm_l_c, n1_adj_519;
    wire [7:0]control_reg_adj_782;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_784;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping_adj_523;
    wire [31:0]read_value_adj_785;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_786;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_558, n3586;
    wire [31:0]n224_adj_789;
    
    wire n14, n27993, n12, n2_adj_591, n10, n32390, n32389, n32388, 
        n32387, n28299, n12031, n12030, bclk;
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    wire [5:0]state_adj_832;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n32386, n7852, n34353, n30658, n6_adj_592, n5, n4_adj_593, 
        n34352, n32369, n15_adj_594, n30940, n32543, n32542, n4_adj_595, 
        n32536, n32534, n30418, n32527, n34351, n28345, n11987, 
        n11981, n11966, n28339, n30520, n32525, n15_adj_596, n32523, 
        n34350, n34349, n2_adj_597, n14_adj_598, n32511, n4_adj_599, 
        n32509, n32508, n2_adj_600, n1_adj_601, n4_adj_602;
    wire [14:0]n66_adj_1126;
    
    wire n4_adj_603, n32503, n4_adj_604, n1_adj_605, n6_adj_606, n16_adj_607, 
        n14_adj_608, n12_adj_609, n10_adj_610, n8, n6_adj_611, n5_adj_612, 
        n4_adj_613, n4_adj_614, n4_adj_615, n1_adj_616, n2_adj_617, 
        n1_adj_618, n2_adj_619, n1_adj_620, n2_adj_621, n1_adj_622, 
        n2_adj_623, n4_adj_624, n1_adj_625, n2_adj_626, n32488, n1_adj_627, 
        n2_adj_628, n1_adj_629, n2_adj_630, n32486, n1_adj_631, n2_adj_632, 
        n1_adj_633, n2_adj_634, n32482, n1_adj_635, n2_adj_636, n1_adj_637, 
        n2_adj_638, n1_adj_639, n2_adj_640, n1_adj_641, n2_adj_642, 
        n1_adj_643, n34348, n30431, n6_adj_644, n29642, n5_adj_645, 
        n32478, n29195, n28337, n30519, n1_adj_646, n14_adj_647, 
        n31642, n31641, n2_adj_648, n32473, n32472, n1_adj_649, 
        n32471, n32469, n32385, n30474, n30454, n30450, n1_adj_650, 
        n30435, n28488;
    wire [12:0]count_adj_843;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    
    wire n30429, n30364, n20291;
    wire [12:0]count_adj_846;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    wire [7:0]n7903;
    
    wire motor_pwm_r_c, n32463, n30316, n30311, n8_adj_658, n32462, 
        n32461, n31041, n15_adj_659, n32, n30743, n30942, n31079, 
        n32454, n32453, n1_adj_660, n2_adj_661, n30839, n34347, 
        n32449, n7902, n29690, n32446, n30831, n32442, n32379, 
        n32441, n30826, n32378, n32375, n14_adj_662, n28214, n2_adj_663, 
        n32438, n32437, n32436, n32435, n8048, n30958, n32430, 
        n30518, n32429, n54, n20418, n30816, n32422, n32420, n32374, 
        n31583, n32416, n12788, n1_adj_664, n2_adj_665, n1_adj_666, 
        n30808, n6674, n32413, n34344, n28401, n32412, n30594, 
        n32411, n30803, n31057, n9_adj_667, n32408, n32407, n32406, 
        n32405, n31050, n988, n1000, n11271;
    
    VHI i2 (.Z(VCC_net));
    PWMPeripheral motor_pwm (.n32478(n32478), .n32488(n32488), .rw(rw), 
            .n34347(n34347), .\read_size[0] (read_size_adj_689[0]), .debug_c_c(debug_c_c), 
            .n30743(n30743), .n34349(n34349), .\databus[0] (databus[0]), 
            .\select[2] (select[2]), .read_value({read_value_adj_688}), 
            .n282(n281[15]), .n34353(n34353), .\databus[6] (databus[6]), 
            .\databus[5] (databus[5]), .\databus[4] (databus[4]), .\databus[3] (databus[3]), 
            .\databus[2] (databus[2]), .\databus[1] (databus[1]), .n32471(n32471), 
            .\register_addr[0] (register_addr[0]), .n34344(n34344), .n64(n64), 
            .\count[0] (count_adj_846[0]), .n32375(n32375), .motor_pwm_r_c(motor_pwm_r_c), 
            .GND_net(GND_net), .n9633(n9633), .n14322(n14322), .\count[1] (count_adj_846[1]), 
            .\count[2] (count_adj_846[2]), .\count[3] (count_adj_846[3]), 
            .\count[4] (count_adj_846[4]), .\count[5] (count_adj_846[5]), 
            .\count[6] (count_adj_846[6]), .\count[7] (count_adj_846[7]), 
            .\count[8] (count_adj_846[8]), .n3589(n3589), .n7893({n7893}), 
            .n7902(n7902), .n10513(n10513), .n14473(n14473), .\count[0]_adj_194 (count_adj_843[0]), 
            .\count[12] (count_adj_843[12]), .\count[11] (count_adj_843[11]), 
            .\count[9] (count_adj_843[9]), .\count[8]_adj_195 (count_adj_843[8]), 
            .\count[6]_adj_196 (count_adj_843[6]), .\count[5]_adj_197 (count_adj_843[5]), 
            .\count[3]_adj_198 (count_adj_843[3]), .\count[2]_adj_199 (count_adj_843[2]), 
            .\count[1]_adj_200 (count_adj_843[1]), .motor_pwm_l_c(motor_pwm_l_c), 
            .n28488(n28488), .n32385(n32385), .n10(n10_adj_610), .n12(n12_adj_609), 
            .\reset_count[6] (reset_count[6]), .n30518(n30518), .\reset_count[4] (reset_count[4]), 
            .\reset_count[5] (reset_count[5]), .n30519(n30519), .n3586(n3586), 
            .n6(n6), .\reset_count[8] (reset_count[8]), .\reset_count[7] (reset_count[7]), 
            .n32430(n32430), .n6_adj_201(n6_adj_611), .n8(n8), .n7912(n7912), 
            .n7906(n7903[5]), .n7905(n7903[6]), .n7908(n7903[3]), .n7910(n7903[1]), 
            .n7909(n7903[2]), .n7911(n7903[0])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(512[16] 522[40])
    LUT4 i24726_4_lut_rep_429 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n34353)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_429.init = 16'h575f;
    LUT4 i1_2_lut_rep_280_3_lut_4_lut (.A(n32482), .B(select[4]), .C(prev_select), 
         .D(n32508), .Z(n32405)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_280_3_lut_4_lut.init = 16'h0004;
    LUT4 i20_2_lut_rep_282_3_lut_4_lut (.A(n32482), .B(select[4]), .C(n34344), 
         .D(n32508), .Z(n32407)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i20_2_lut_rep_282_3_lut_4_lut.init = 16'h0040;
    LUT4 i20_2_lut_rep_281_3_lut_4_lut (.A(n32482), .B(select[4]), .C(rw), 
         .D(n30454), .Z(n32406)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i20_2_lut_rep_281_3_lut_4_lut.init = 16'h4000;
    LUT4 n9396_c_bdd_4_lut (.A(n9396_c), .B(state_adj_832[1]), .C(rdata[1]), 
         .D(bclk), .Z(n31641)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam n9396_c_bdd_4_lut.init = 16'hb8f0;
    LUT4 i1_2_lut_rep_291_3_lut_4_lut (.A(n32482), .B(select[4]), .C(prev_select_adj_558), 
         .D(n30454), .Z(n32416)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_291_3_lut_4_lut.init = 16'h0400;
    LUT4 i20_2_lut_rep_283_3_lut_4_lut (.A(n32482), .B(select[4]), .C(rw), 
         .D(n32534), .Z(n32408)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i20_2_lut_rep_283_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_297_3_lut_4_lut (.A(n32482), .B(select[4]), .C(prev_select_adj_518), 
         .D(n32534), .Z(n32422)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_297_3_lut_4_lut.init = 16'h0004;
    PFUMX LessThan_1437_i18 (.BLUT(n14), .ALUT(n16), .C0(n30839), .Z(n3589));
    PFUMX LessThan_1434_i18 (.BLUT(n14_adj_608), .ALUT(n16_adj_607), .C0(n30816), 
          .Z(n3586));
    PFUMX i22 (.BLUT(n15_adj_594), .ALUT(n30934), .C0(state_adj_832[0]), 
          .Z(n29195));
    LUT4 LessThan_1434_i13_2_lut_rep_278 (.A(n7903[6]), .B(count_adj_843[6]), 
         .Z(n32403)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i13_2_lut_rep_278.init = 16'h6666;
    LUT4 LessThan_1434_i10_3_lut_3_lut (.A(n7903[6]), .B(count_adj_843[6]), 
         .C(count_adj_843[5]), .Z(n10_adj_610)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1434_i11_2_lut_rep_279 (.A(n7903[5]), .B(count_adj_843[5]), 
         .Z(n32404)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i11_2_lut_rep_279.init = 16'h6666;
    LUT4 i24450_2_lut_3_lut_4_lut (.A(n7903[5]), .B(count_adj_843[5]), .C(count_adj_843[6]), 
         .D(n7903[6]), .Z(n30808)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24450_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 Select_3599_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[17]), 
         .D(rw), .Z(n1_adj_633)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3599_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3597_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[18]), 
         .D(rw), .Z(n1_adj_637)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3597_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i14030_2_lut_2_lut (.A(n34347), .B(databus[0]), .Z(n571[0])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14030_2_lut_2_lut.init = 16'h4444;
    LUT4 n32525_bdd_4_lut (.A(n32525), .B(n32527), .C(register_addr[1]), 
         .D(register_addr[0]), .Z(n30450)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n32525_bdd_4_lut.init = 16'h0010;
    LUT4 Select_3595_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[19]), 
         .D(rw), .Z(n2_adj_632)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3595_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3599_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[17]), 
         .D(rw), .Z(n2_adj_634)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3599_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3597_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[18]), 
         .D(rw), .Z(n2_adj_638)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3597_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3601_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[16]), 
         .D(rw), .Z(n2_adj_642)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3601_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3603_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[15]), 
         .D(rw), .Z(n2_adj_640)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3603_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3605_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[14]), 
         .D(rw), .Z(n2_adj_630)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3605_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_2_lut_rep_311_3_lut_4_lut (.A(n32543), .B(n32542), .C(state_adj_832[5]), 
         .D(state_adj_832[0]), .Z(n32436)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i2_2_lut_rep_311_3_lut_4_lut.init = 16'h0010;
    LUT4 Select_3607_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[13]), 
         .D(rw), .Z(n2_adj_628)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3607_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3609_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[12]), 
         .D(rw), .Z(n2_adj_626)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3609_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_4_lut (.A(state_adj_832[5]), .B(state_adj_832[1]), .C(n183), 
         .D(n32), .Z(n15_adj_594)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_4_lut.init = 16'h4505;
    LUT4 i24667_2_lut (.A(bclk), .B(state_adj_832[1]), .Z(n30934)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i24667_2_lut.init = 16'h9999;
    LUT4 Select_3611_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[11]), 
         .D(rw), .Z(n2_adj_621)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3611_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3613_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[10]), 
         .D(rw), .Z(n2_adj_617)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3613_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3615_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[9]), 
         .D(rw), .Z(n2_adj_623)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3615_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3617_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[8]), 
         .D(rw), .Z(n2_adj_619)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3617_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3571_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[31]), 
         .D(rw), .Z(n2_adj_600)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3571_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3577_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[28]), 
         .D(rw), .Z(n2_adj_442)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3577_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3573_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[30]), 
         .D(rw), .Z(n2_adj_597)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3573_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3575_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[29]), 
         .D(rw), .Z(n2_adj_663)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3575_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3579_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[27]), 
         .D(rw), .Z(n2)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3579_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3581_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[26]), 
         .D(rw), .Z(n2_adj_394)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3581_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3583_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[25]), 
         .D(rw), .Z(n2_adj_648)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3583_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3585_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[24]), 
         .D(rw), .Z(n2_adj_661)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3585_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3587_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[23]), 
         .D(rw), .Z(n2_adj_396)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3587_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3589_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[22]), 
         .D(rw), .Z(n2_adj_665)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3589_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3591_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[21]), 
         .D(rw), .Z(n2_adj_591)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3591_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3593_i2_2_lut_3_lut_4_lut (.A(n32534), .B(n32469), .C(read_value_adj_745[20]), 
         .D(rw), .Z(n2_adj_636)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3593_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_271_3_lut_4_lut (.A(n32534), .B(n32469), .C(rw), 
         .D(prev_select_adj_518), .Z(n32396)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_271_3_lut_4_lut.init = 16'h0004;
    LUT4 i24726_4_lut_rep_423 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n34347)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_423.init = 16'h575f;
    LUT4 i2_3_lut_rep_275_4_lut_4_lut (.A(n34347), .B(n30311), .C(prev_select_adj_518), 
         .D(n32449), .Z(n32400)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_275_4_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n34347), .B(register_addr[1]), .C(n30311), 
         .D(n32422), .Z(n30316)) /* synthesis lut_function=(A (B)+!A (B (C+!(D)))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'hc8cc;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n34347), .B(prev_select_adj_518), 
         .C(n32469), .D(n32534), .Z(n11981)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_471 (.A(n34347), .B(prev_select), 
         .C(n32469), .D(n32508), .Z(n11966)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_471.init = 16'h0010;
    LUT4 i13958_2_lut_2_lut (.A(n34347), .B(n6674), .Z(n241)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i13958_2_lut_2_lut.init = 16'h4444;
    LUT4 i13999_2_lut_2_lut (.A(n34347), .B(databus[7]), .Z(n281[15])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i13999_2_lut_2_lut.init = 16'h4444;
    LUT4 i24750_4_lut_4_lut (.A(n32472), .B(n4_adj_479), .C(n9_adj_667), 
         .D(n1286[14]), .Z(n12098)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i24750_4_lut_4_lut.init = 16'h2a00;
    LUT4 i3_4_lut_4_lut (.A(n32472), .B(n32536), .C(n1286[8]), .D(n1286[0]), 
         .Z(n12788)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i3_4_lut_4_lut.init = 16'hfffd;
    LUT4 i24726_4_lut_rep_424 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n34348)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_424.init = 16'h575f;
    LUT4 i1_2_lut_rep_383 (.A(register_addr[4]), .B(register_addr[5]), .Z(n32508)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i1_2_lut_rep_383.init = 16'heeee;
    LUT4 i24252_2_lut_rep_337_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(register_addr[0]), .D(n32509), .Z(n32462)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i24252_2_lut_rep_337_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_rep_329_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(n32527), .D(n32509), .Z(n32454)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i2_2_lut_rep_329_3_lut_4_lut.init = 16'hfffe;
    LUT4 LessThan_1434_i17_2_lut_rep_261 (.A(n7912), .B(count_adj_843[8]), 
         .Z(n32386)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i17_2_lut_rep_261.init = 16'h6666;
    FD1P3AX reset_count_2172_2173__i1 (.D(n66_adj_1126[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i1.GSR = "ENABLED";
    LUT4 LessThan_1434_i16_3_lut_3_lut (.A(n7912), .B(count_adj_843[8]), 
         .C(n8), .Z(n16_adj_607)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24726_4_lut_rep_425 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n34349)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_425.init = 16'h575f;
    LUT4 Select_3595_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[19]), 
         .D(rw), .Z(n1_adj_631)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3595_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3603_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[15]), 
         .D(rw), .Z(n1_adj_639)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3603_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3605_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[14]), 
         .D(rw), .Z(n1_adj_629)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3605_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 n227_bdd_4_lut (.A(n9396_c), .B(state_adj_832[1]), .C(rdata[0]), 
         .D(bclk), .Z(n31582)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam n227_bdd_4_lut.init = 16'he2f0;
    LUT4 i24726_4_lut_rep_426 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n34350)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_426.init = 16'h575f;
    LUT4 Select_3607_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[13]), 
         .D(rw), .Z(n1_adj_627)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3607_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1437_i15_2_lut_rep_264 (.A(n7893[7]), .B(count_adj_846[7]), 
         .Z(n32389)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i15_2_lut_rep_264.init = 16'h6666;
    LUT4 LessThan_1437_i12_3_lut_3_lut (.A(n7893[7]), .B(count_adj_846[7]), 
         .C(n10), .Z(n12)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1437_i17_2_lut_rep_265 (.A(n7902), .B(count_adj_846[8]), 
         .Z(n32390)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i17_2_lut_rep_265.init = 16'h6666;
    LUT4 LessThan_1437_i16_3_lut_3_lut (.A(n7902), .B(count_adj_846[8]), 
         .C(n8_adj_658), .Z(n16)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_rep_321_4_lut (.A(select[4]), .B(n32482), .C(n30283), 
         .D(prev_select_adj_478), .Z(n32446)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i1_2_lut_rep_321_4_lut.init = 16'h0020;
    LUT4 i20_2_lut_4_lut (.A(select[4]), .B(n32482), .C(n30283), .D(rw), 
         .Z(n52)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i20_2_lut_4_lut.init = 16'h2000;
    LUT4 i1_4_lut_adj_472 (.A(n19896), .B(reset_count[11]), .C(reset_count[8]), 
         .D(n27993), .Z(n30429)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_472.init = 16'h8880;
    LUT4 i2_3_lut (.A(reset_count[7]), .B(reset_count[5]), .C(reset_count[6]), 
         .Z(n27993)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i24726_4_lut_rep_338 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n32463)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_338.init = 16'h575f;
    LUT4 i24726_4_lut_rep_427 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n34351)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_427.init = 16'h575f;
    LUT4 Select_3609_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[12]), 
         .D(n34344), .Z(n1_adj_625)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3609_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24726_4_lut_rep_428 (.A(reset_count[14]), .B(n30519), .C(n29642), 
         .D(n19896), .Z(n34352)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24726_4_lut_rep_428.init = 16'h575f;
    LUT4 Select_3611_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[11]), 
         .D(n34344), .Z(n1_adj_620)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3611_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    IB n9396_pad (.I(uart_rx), .O(n9396_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    OB debug_pad_0 (.I(n9396_c), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_1 (.I(n9395), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_6 (.I(n34347), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB motor_pwm_r_pad (.I(motor_pwm_r_c), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    LUT4 Select_3613_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[10]), 
         .D(n34344), .Z(n1_adj_616)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3613_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    OB expansion5_pad (.I(GND_net), .O(expansion5));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    OB expansion4_pad (.I(GND_net), .O(expansion4));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    OB expansion3_pad (.I(GND_net), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    OB expansion2_pad (.I(GND_net), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion1_pad (.I(GND_net), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    LUT4 Select_3615_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[9]), 
         .D(rw), .Z(n1_adj_622)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3615_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB uart_tx_pad (.I(n9395), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    LUT4 Select_3617_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[8]), 
         .D(rw), .Z(n1_adj_618)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3617_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_adj_473 (.A(reset_count[12]), .B(reset_count[13]), .C(reset_count[11]), 
         .Z(n29642)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[17:42])
    defparam i2_3_lut_adj_473.init = 16'hfefe;
    LUT4 i1_2_lut_rep_417 (.A(state_adj_832[1]), .B(state_adj_832[4]), .Z(n32542)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_rep_417.init = 16'heeee;
    LUT4 i1_2_lut_rep_336_3_lut_4_lut (.A(state_adj_832[1]), .B(state_adj_832[4]), 
         .C(state_adj_832[0]), .D(n32543), .Z(n32461)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_rep_336_3_lut_4_lut.init = 16'hfffe;
    LUT4 Select_3571_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[31]), 
         .D(rw), .Z(n1_adj_601)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3571_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state_adj_832[1]), .B(state_adj_832[4]), 
         .C(n9396_c), .D(n32543), .Z(n183)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_418 (.A(state_adj_832[2]), .B(state_adj_832[3]), .Z(n32543)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_rep_418.init = 16'heeee;
    LUT4 n31641_bdd_3_lut_4_lut (.A(state_adj_832[2]), .B(state_adj_832[3]), 
         .C(rdata[1]), .D(n31641), .Z(n31642)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam n31641_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n31582_bdd_3_lut_4_lut (.A(state_adj_832[2]), .B(state_adj_832[3]), 
         .C(rdata[0]), .D(n31582), .Z(n31583)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam n31582_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24661_4_lut (.A(n4), .B(n12), .C(n32389), .D(n30831), .Z(n14)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24661_4_lut.init = 16'hcacc;
    LUT4 LessThan_1437_i4_4_lut (.A(count_adj_846[0]), .B(count_adj_846[1]), 
         .C(n7893[1]), .D(n7893[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i4_4_lut.init = 16'h8ecf;
    LUT4 i24811_4_lut (.A(n32390), .B(n32389), .C(n32411), .D(n30826), 
         .Z(n30839)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24811_4_lut.init = 16'habaa;
    LUT4 i24468_4_lut (.A(n32412), .B(n32438), .C(n32437), .D(n5_adj_645), 
         .Z(n30826)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24468_4_lut.init = 16'h5554;
    LUT4 LessThan_1437_i5_2_lut (.A(n7893[2]), .B(count_adj_846[2]), .Z(n5_adj_645)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i5_2_lut.init = 16'h6666;
    FD1P3AX reset_count_2172_2173__i2 (.D(n66_adj_1126[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i2.GSR = "ENABLED";
    LUT4 i3_4_lut_rep_244 (.A(n54), .B(n6_adj_439), .C(n1000), .D(n4_adj_595), 
         .Z(n32369)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+!(D))+!B))) */ ;
    defparam i3_4_lut_rep_244.init = 16'h0c08;
    LUT4 i8680_2_lut_3_lut (.A(n54), .B(n6_adj_439), .C(n1000), .Z(n14446)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i8680_2_lut_3_lut.init = 16'h0808;
    LUT4 Select_3577_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[28]), 
         .D(rw), .Z(n1_adj_649)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3577_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3573_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[30]), 
         .D(n34344), .Z(n1_adj_646)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3573_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3575_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[29]), 
         .D(n34344), .Z(n1_adj_519)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3575_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3579_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[27]), 
         .D(n34344), .Z(n1)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3579_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    GSR GSR_INST (.GSR(VCC_net));
    FD1P3AX reset_count_2172_2173__i3 (.D(n66_adj_1126[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i4 (.D(n66_adj_1126[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i5 (.D(n66_adj_1126[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i6 (.D(n66_adj_1126[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i7 (.D(n66_adj_1126[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i8 (.D(n66_adj_1126[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i9 (.D(n66_adj_1126[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i10 (.D(n66_adj_1126[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i11 (.D(n66_adj_1126[10]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i12 (.D(n66_adj_1126[11]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i13 (.D(n66_adj_1126[12]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i14 (.D(n66_adj_1126[13]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i15 (.D(n66_adj_1126[14]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i15.GSR = "ENABLED";
    LUT4 Select_3581_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[26]), 
         .D(n34344), .Z(n1_adj_395)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3581_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1437_i13_2_lut_rep_286 (.A(n7893[6]), .B(count_adj_846[6]), 
         .Z(n32411)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i13_2_lut_rep_286.init = 16'h6666;
    LUT4 i24757_4_lut (.A(count_adj_843[9]), .B(count_adj_843[11]), .C(count_adj_843[12]), 
         .D(n6), .Z(n28488)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24757_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut (.A(n32395), .B(n30450), .C(n34347), .Z(n12224)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 Select_3583_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[25]), 
         .D(n34344), .Z(n1_adj_650)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3583_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(register_addr[4]), .B(register_addr[5]), .Z(n30283)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 LessThan_1437_i10_3_lut_3_lut (.A(n7893[6]), .B(count_adj_846[6]), 
         .C(count_adj_846[5]), .Z(n10)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 Select_3585_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[24]), 
         .D(n34344), .Z(n1_adj_660)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3585_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    VLO i1 (.Z(GND_net));
    LUT4 Select_3587_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[23]), 
         .D(n34344), .Z(n1_adj_664)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3587_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24695_4_lut (.A(n30520), .B(reset_count[14]), .C(n29642), .D(n19896), 
         .Z(n30)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i24695_4_lut.init = 16'h373f;
    LUT4 i1_4_lut_adj_474 (.A(n20418), .B(n30518), .C(reset_count[6]), 
         .D(reset_count[5]), .Z(n30520)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[7:30])
    defparam i1_4_lut_adj_474.init = 16'hfcec;
    LUT4 i14680_4_lut (.A(reset_count[0]), .B(reset_count[4]), .C(n6_adj_393), 
         .D(reset_count[3]), .Z(n20418)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i14680_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(reset_count[1]), .B(reset_count[2]), .Z(n6_adj_393)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i24659_4_lut (.A(n4_adj_613), .B(n12_adj_609), .C(n32385), .D(n30808), 
         .Z(n14_adj_608)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24659_4_lut.init = 16'hcacc;
    LUT4 LessThan_1434_i7_2_lut_rep_304 (.A(n7903[3]), .B(count_adj_843[3]), 
         .Z(n32429)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i7_2_lut_rep_304.init = 16'h6666;
    LUT4 LessThan_1434_i6_3_lut_3_lut (.A(n7903[3]), .B(count_adj_843[3]), 
         .C(count_adj_843[2]), .Z(n6_adj_611)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1437_i7_2_lut_rep_312 (.A(n7893[3]), .B(count_adj_846[3]), 
         .Z(n32437)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i7_2_lut_rep_312.init = 16'h6666;
    LUT4 Select_3589_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[22]), 
         .D(n34344), .Z(n1_adj_666)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3589_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3591_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[21]), 
         .D(n34344), .Z(n1_adj_643)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3591_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1437_i6_3_lut_3_lut (.A(n7893[3]), .B(count_adj_846[3]), 
         .C(count_adj_846[2]), .Z(n6_adj_644)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i2_3_lut_rep_263_4_lut_4_lut (.A(n34347), .B(n32454), .C(prev_select), 
         .D(n32435), .Z(n32388)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_rep_263_4_lut_4_lut.init = 16'h0400;
    LUT4 Select_3593_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[20]), 
         .D(n34344), .Z(n1_adj_635)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3593_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1434_i4_4_lut (.A(count_adj_843[0]), .B(count_adj_843[1]), 
         .C(n7903[1]), .D(n7903[0]), .Z(n4_adj_613)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i4_4_lut.init = 16'h8ecf;
    LUT4 i1_2_lut_4_lut_4_lut_adj_475 (.A(n34347), .B(register_addr[1]), 
         .C(n32454), .D(n32405), .Z(n30364)) /* synthesis lut_function=(A (B)+!A !((C (D))+!B)) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_475.init = 16'h8ccc;
    LUT4 i14005_2_lut_2_lut (.A(n34347), .B(databus[4]), .Z(n580[4])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14005_2_lut_2_lut.init = 16'h4444;
    LUT4 LessThan_1437_i9_2_lut_rep_313 (.A(n7893[4]), .B(count_adj_846[4]), 
         .Z(n32438)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i9_2_lut_rep_313.init = 16'h6666;
    LUT4 i1_3_lut_rep_270_4_lut_4_lut (.A(n32469), .B(n30454), .C(n34344), 
         .D(prev_select_adj_558), .Z(n32395)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_270_4_lut_4_lut.init = 16'h0008;
    LUT4 LessThan_1437_i8_3_lut_3_lut (.A(n7893[4]), .B(count_adj_846[4]), 
         .C(n6_adj_644), .Z(n8_adj_658)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24837_4_lut (.A(n32386), .B(n32385), .C(n32403), .D(n30803), 
         .Z(n30816)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24837_4_lut.init = 16'habaa;
    LUT4 i24445_4_lut (.A(n32404), .B(n32430), .C(n32429), .D(n5_adj_612), 
         .Z(n30803)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24445_4_lut.init = 16'h5554;
    LUT4 LessThan_1437_i11_2_lut_rep_287 (.A(n7893[5]), .B(count_adj_846[5]), 
         .Z(n32412)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i11_2_lut_rep_287.init = 16'h6666;
    LUT4 i24473_2_lut_3_lut_4_lut (.A(n7893[5]), .B(count_adj_846[5]), .C(count_adj_846[6]), 
         .D(n7893[6]), .Z(n30831)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24473_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 LessThan_1434_i5_2_lut (.A(n7903[2]), .B(count_adj_843[2]), .Z(n5_adj_612)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i5_2_lut.init = 16'h6666;
    LUT4 i14127_2_lut_2_lut (.A(n34347), .B(databus[2]), .Z(n580[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14127_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_262_3_lut_4_lut (.A(n32508), .B(n32469), .C(rw), 
         .D(prev_select), .Z(n32387)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_262_3_lut_4_lut.init = 16'h0004;
    LUT4 Select_3621_i4_2_lut_3_lut_4_lut (.A(n32508), .B(n32469), .C(read_value_adj_693[4]), 
         .D(n34344), .Z(n4_adj_614)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3621_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3622_i4_2_lut_3_lut_4_lut (.A(n32508), .B(n32469), .C(read_value_adj_693[3]), 
         .D(n34344), .Z(n4_adj_604)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3622_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3623_i4_2_lut_3_lut_4_lut (.A(n32508), .B(n32469), .C(read_value_adj_693[2]), 
         .D(n34344), .Z(n4_adj_603)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3623_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3625_i4_2_lut_3_lut_4_lut (.A(n32508), .B(n32469), .C(read_value_adj_693[0]), 
         .D(rw), .Z(n4_adj_602)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3625_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    GlobalControlPeripheral global_control (.read_value({read_value[31:2], 
            Open_0, read_value[0]}), .debug_c_c(debug_c_c), .n32413(n32413), 
            .register_addr({register_addr}), .n32486(n32486), .n8048(n8048), 
            .n11753(n11753), .n30418(n30418), .read_size({read_size}), 
            .n302(n302), .\register[2] ({Open_1, Open_2, Open_3, Open_4, 
            Open_5, Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, 
            Open_12, Open_13, Open_14, Open_15, Open_16, Open_17, 
            Open_18, Open_19, Open_20, Open_21, Open_22, Open_23, 
            Open_24, Open_25, Open_26, Open_27, Open_28, Open_29, 
            Open_30, Open_31, \register[2] [0]}), .n34348(n34348), .\select[1] (select[1]), 
            .\select[4] (select[4]), .n32527(n32527), .n32469(n32469), 
            .n32454(n32454), .n34350(n34350), .n34349(n34349), .\register[2][3] (\register[2] [3]), 
            .n28386(n28386), .n32453(n32453), .n32463(n32463), .n15(n15_adj_596), 
            .n32462(n32462), .n4(n4_adj_593), .n10513(n10513), .n14473(n14473), 
            .signal_light_c(signal_light_c), .n9633(n9633), .n14322(n14322), 
            .\control_reg[7] (control_reg[7]), .n28360(n28360), .n18(n18), 
            .\control_reg[7]_adj_188 (control_reg_adj_782[7]), .n28299(n28299), 
            .stepping(stepping_adj_523), .\control_reg[7]_adj_189 (control_reg_adj_702[7]), 
            .n28401(n28401), .stepping_adj_190(stepping), .\control_reg[7]_adj_191 (control_reg_adj_742[7]), 
            .n28214(n28214), .stepping_adj_192(stepping_adj_483), .rw(rw), 
            .n32503(n32503), .n6(n6_adj_606), .n32478(n32478), .n11645(n11645), 
            .\databus[1] (databus[1]), .n34347(n34347), .n32525(n32525), 
            .xbee_pause_c(xbee_pause_c), .n20291(n20291), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(495[45] 505[74])
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.n34344(n34344), .n32422(n32422), 
            .\register_addr[5] (register_addr[5]), .n30431(n30431), .read_value({read_value_adj_745}), 
            .debug_c_c(debug_c_c), .n11981(n11981), .n32400(n32400), .\register_addr[1] (register_addr[1]), 
            .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_Z_nFault_c(Stepper_Z_nFault_c), 
            .n34349(n34349), .\read_size[0] (read_size_adj_746[0]), .n30658(n30658), 
            .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n579(n571[0]), .prev_select(prev_select_adj_518), 
            .n32449(n32449), .n32534(n32534), .n32442(n32442), .rw(rw), 
            .n34347(n34347), .n32396(n32396), .n7852(n7852), .n34350(n34350), 
            .databus({databus}), .n608(n580[4]), .n610(n580[2]), .\control_reg[7] (control_reg_adj_742[7]), 
            .Stepper_Z_En_c(Stepper_Z_En_c), .n34351(n34351), .Stepper_Z_Dir_c(Stepper_Z_Dir_c), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), 
            .\read_size[2] (read_size_adj_746[2]), .n29690(n29690), .\steps_reg[5] (steps_reg_adj_744[5]), 
            .\steps_reg[3] (steps_reg_adj_744[3]), .n34352(n34352), .n14(n14_adj_598), 
            .\register_addr[0] (register_addr[0]), .n15(n15_adj_440), .stepping(stepping_adj_483), 
            .n30316(n30316), .n32473(n32473), .n32525(n32525), .n32395(n32395), 
            .n20528(n20528), .limit_c_2(limit_c_2), .n28214(n28214), .Stepper_Z_Step_c(Stepper_Z_Step_c), 
            .n32463(n32463)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(589[25] 602[45])
    LUT4 Select_3618_i4_2_lut_3_lut_4_lut (.A(n32508), .B(n32469), .C(read_value_adj_693[7]), 
         .D(rw), .Z(n4_adj_624)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3618_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3619_i4_2_lut_3_lut_4_lut (.A(n32508), .B(n32469), .C(read_value_adj_693[6]), 
         .D(rw), .Z(n4_adj_599)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3619_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3620_i4_2_lut_3_lut_4_lut (.A(n32508), .B(n32469), .C(read_value_adj_693[5]), 
         .D(rw), .Z(n4_adj_615)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3620_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.register_addr({register_addr}), 
            .read_value({read_value_adj_785}), .debug_c_c(debug_c_c), .n12620(n12620), 
            .GND_net(GND_net), .n34350(n34350), .n3181({n3181}), .VCC_net(VCC_net), 
            .Stepper_A_nFault_c(Stepper_A_nFault_c), .\read_size[0] (read_size_adj_786[0]), 
            .n30435(n30435), .n32527(n32527), .n32525(n32525), .n30311(n30311), 
            .Stepper_A_M0_c_0(Stepper_A_M0_c_0), .n20528(n20528), .n579(n571[0]), 
            .n12224(n12224), .prev_select(prev_select_adj_558), .n32441(n32441), 
            .n32379(n32379), .n34348(n34348), .\databus[31] (databus[31]), 
            .\databus[28] (databus[28]), .n34349(n34349), .\databus[13] (databus[13]), 
            .\databus[11] (databus[11]), .\databus[10] (databus[10]), .\databus[9] (databus[9]), 
            .\databus[7] (databus[7]), .\databus[6] (databus[6]), .\databus[5] (databus[5]), 
            .n610(n580[2]), .\control_reg[7] (control_reg_adj_782[7]), .Stepper_A_En_c(Stepper_A_En_c), 
            .Stepper_A_Dir_c(Stepper_A_Dir_c), .\databus[4] (databus[4]), 
            .\databus[3] (databus[3]), .Stepper_A_M2_c_2(Stepper_A_M2_c_2), 
            .Stepper_A_M1_c_1(Stepper_A_M1_c_1), .\databus[1] (databus[1]), 
            .\read_size[2] (read_size_adj_786[2]), .n30363(n30363), .n32396(n32396), 
            .n7852(n7852), .n34351(n34351), .n34352(n34352), .\steps_reg[5] (steps_reg_adj_784[5]), 
            .\steps_reg[3] (steps_reg_adj_784[3]), .n32442(n32442), .n32508(n32508), 
            .n32509(n32509), .n32471(n32471), .n14(n14_adj_662), .n15(n15_adj_659), 
            .n224({n224_adj_789}), .n32482(n32482), .\register[2][0] (\register[2] [0]), 
            .n15_adj_187(n15_adj_596), .\register[2][3] (\register[2] [3]), 
            .n4(n4_adj_593), .n32488(n32488), .n32473(n32473), .stepping(stepping_adj_523), 
            .n34347(n34347), .\databus[8] (databus[8]), .\databus[12] (databus[12]), 
            .\databus[14] (databus[14]), .\databus[15] (databus[15]), .\databus[16] (databus[16]), 
            .\databus[17] (databus[17]), .\databus[18] (databus[18]), .\databus[19] (databus[19]), 
            .\databus[20] (databus[20]), .\databus[21] (databus[21]), .\databus[22] (databus[22]), 
            .\databus[23] (databus[23]), .\databus[24] (databus[24]), .\databus[25] (databus[25]), 
            .\databus[26] (databus[26]), .\databus[27] (databus[27]), .\databus[29] (databus[29]), 
            .\databus[30] (databus[30]), .limit_c_3(limit_c_3), .n32416(n32416), 
            .n30454(n30454), .rw(rw), .n28299(n28299), .Stepper_A_Step_c(Stepper_A_Step_c), 
            .n32463(n32463)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(604[25] 617[45])
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_476 (.A(n34347), .B(prev_select_adj_558), 
         .C(n30454), .D(n32469), .Z(n12620)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_476.init = 16'h1000;
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.\register_addr[1] (register_addr[1]), 
            .databus({databus}), .n3363(n3363), .debug_c_c(debug_c_c), 
            .n34349(n34349), .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .\read_size[0] (read_size_adj_706[0]), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), 
            .n579(n571[0]), .\register_addr[0] (register_addr[0]), .n12434(n12434), 
            .prev_select(prev_select_adj_478), .n32523(n32523), .n32509(n32509), 
            .n32527(n32527), .n32525(n32525), .n30283(n30283), .\select[4] (select[4]), 
            .n32508(n32508), .n32435(n32435), .n30454(n30454), .n32441(n32441), 
            .n32534(n32534), .n32449(n32449), .read_value({read_value_adj_705}), 
            .n34348(n34348), .n34351(n34351), .n34350(n34350), .n34352(n34352), 
            .\control_reg[7] (control_reg_adj_702[7]), .Stepper_Y_En_c(Stepper_Y_En_c), 
            .Stepper_Y_Dir_c(Stepper_Y_Dir_c), .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), 
            .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), .\read_size[2] (read_size_adj_706[2]), 
            .n30474(n30474), .n34353(n34353), .\steps_reg[5] (steps_reg_adj_704[5]), 
            .\steps_reg[3] (steps_reg_adj_704[3]), .n34344(n34344), .n32420(n32420), 
            .n34347(n34347), .n14(n14_adj_647), .n15(n15), .limit_c_1(limit_c_1), 
            .stepping(stepping), .\register_addr[5] (register_addr[5]), 
            .\register_addr[4] (register_addr[4]), .n32442(n32442), .rw(rw), 
            .n32446(n32446), .n30450(n30450), .Stepper_Y_Step_c(Stepper_Y_Step_c), 
            .n28401(n28401), .n32463(n32463)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(574[25] 587[45])
    LUT4 Select_3624_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[1]), 
         .D(rw), .Z(n1_adj_605)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3624_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    RCPeripheral rc_receiver (.\register_addr[0] (register_addr[0]), .databus_out({databus_out}), 
            .n2(n2_adj_628), .rw(rw), .databus({databus}), .\read_value[13] (read_value[13]), 
            .n1(n1_adj_627), .n32503(n32503), .\read_value[13]_adj_43 (read_value_adj_693[13]), 
            .read_value({read_value_adj_705}), .n32407(n32407), .n52(n52), 
            .n2_adj_45(n2_adj_626), .\read_value[12]_adj_46 (read_value[12]), 
            .n1_adj_47(n1_adj_625), .\read_value[12]_adj_48 (read_value_adj_693[12]), 
            .\register_addr[2] (register_addr[2]), .\register_addr[1] (register_addr[1]), 
            .n2_adj_49(n2_adj_632), .\select[7] (select[7]), .n32527(n32527), 
            .n32509(n32509), .n30454(n30454), .n30363(n30363), .n32523(n32523), 
            .n30474(n30474), .n32534(n32534), .n30658(n30658), .n29690(n29690), 
            .n30435(n30435), .n2_adj_50(n2_adj_621), .\read_value[11]_adj_51 (read_value[11]), 
            .n1_adj_52(n1_adj_620), .\read_value[11]_adj_53 (read_value_adj_693[11]), 
            .n2_adj_54(n2_adj_617), .\read_value[10]_adj_55 (read_value[10]), 
            .n1_adj_56(n1_adj_616), .\read_value[10]_adj_57 (read_value_adj_693[10]), 
            .\register_addr[4] (register_addr[4]), .n2_adj_58(n2_adj_638), 
            .\read_value[18]_adj_59 (read_value[18]), .n1_adj_60(n1_adj_637), 
            .\read_value[18]_adj_61 (read_value_adj_693[18]), .\read_size[0] (read_size_adj_694[0]), 
            .\read_size[0]_adj_62 (read_size_adj_746[0]), .\register_addr[5] (register_addr[5]), 
            .\read_size[0]_adj_63 (read_size_adj_706[0]), .\read_size[0]_adj_64 (read_size_adj_786[0]), 
            .read_size({read_size}), .\select[1] (select[1]), .n32511(n32511), 
            .\sendcount[1] (sendcount[1]), .n11271(n11271), .n2_adj_66(n2_adj_623), 
            .\read_value[19]_adj_67 (read_value[19]), .n1_adj_68(n1_adj_631), 
            .\read_value[9]_adj_69 (read_value[9]), .n1_adj_70(n1_adj_622), 
            .n2_adj_71(n2_adj_648), .\read_value[25]_adj_72 (read_value[25]), 
            .n1_adj_73(n1_adj_650), .n2_adj_74(n2_adj_636), .\read_value[9]_adj_75 (read_value_adj_693[9]), 
            .\read_value[19]_adj_76 (read_value_adj_693[19]), .n2_adj_77(n2_adj_634), 
            .\read_value[17]_adj_78 (read_value[17]), .n1_adj_79(n1_adj_633), 
            .\read_value[17]_adj_80 (read_value_adj_693[17]), .n2_adj_81(n2_adj_642), 
            .\read_value[20]_adj_82 (read_value[20]), .n1_adj_83(n1_adj_635), 
            .\read_value[16]_adj_84 (read_value[16]), .n1_adj_85(n1_adj_641), 
            .\read_value[16]_adj_86 (read_value_adj_693[16]), .\read_value[25]_adj_87 (read_value_adj_693[25]), 
            .n32486(n32486), .\register_addr[3] (register_addr[3]), .n30594(n30594), 
            .n2_adj_88(n2_adj_640), .\read_value[15]_adj_89 (read_value[15]), 
            .n1_adj_90(n1_adj_639), .n2_adj_91(n2_adj_619), .\read_value[15]_adj_92 (read_value_adj_693[15]), 
            .\read_value[8]_adj_93 (read_value[8]), .n1_adj_94(n1_adj_618), 
            .n2_adj_95(n2_adj_630), .\read_value[14]_adj_96 (read_value[14]), 
            .n1_adj_97(n1_adj_629), .n2_adj_98(n2_adj_597), .\read_value[14]_adj_99 (read_value_adj_693[14]), 
            .\read_value[30]_adj_100 (read_value[30]), .n1_adj_101(n1_adj_646), 
            .n32416(n32416), .n30450(n30450), .n32379(n32379), .\read_value[8]_adj_102 (read_value_adj_693[8]), 
            .n2_adj_103(n2_adj_661), .\select[2] (select[2]), .\read_size[0]_adj_104 (read_size_adj_689[0]), 
            .n5(n5), .n32469(n32469), .n6(n6_adj_592), .\reg_size[2] (reg_size[2]), 
            .\read_value[24]_adj_105 (read_value[24]), .n1_adj_106(n1_adj_660), 
            .\read_value[24]_adj_107 (read_value_adj_693[24]), .\read_value[20]_adj_108 (read_value_adj_693[20]), 
            .n4(n4_adj_624), .\read_value[7]_adj_109 (read_value_adj_785[7]), 
            .n32406(n32406), .\read_value[7]_adj_110 (read_value_adj_745[7]), 
            .\read_value[7]_adj_111 (read_value[7]), .n32408(n32408), .n34344(n34344), 
            .read_value_adj_186({read_value_adj_688}), .n64(n64), .n4_adj_120(n4_adj_599), 
            .\read_value[6]_adj_121 (read_value_adj_785[6]), .\read_value[6]_adj_122 (read_value_adj_745[6]), 
            .\read_value[6]_adj_123 (read_value[6]), .\read_value[30]_adj_124 (read_value_adj_693[30]), 
            .n2_adj_125(n2_adj_396), .\read_value[23]_adj_126 (read_value[23]), 
            .n1_adj_127(n1_adj_664), .n4_adj_128(n4_adj_615), .\read_value[23]_adj_129 (read_value_adj_693[23]), 
            .\read_value[5]_adj_130 (read_value_adj_785[5]), .\read_value[5]_adj_131 (read_value_adj_745[5]), 
            .\read_value[5]_adj_132 (read_value[5]), .n4_adj_133(n4_adj_614), 
            .\read_value[4]_adj_134 (read_value_adj_785[4]), .\read_value[4]_adj_135 (read_value_adj_745[4]), 
            .\read_value[4]_adj_136 (read_value[4]), .n2_adj_137(n2_adj_665), 
            .\read_value[22]_adj_138 (read_value[22]), .n1_adj_139(n1_adj_666), 
            .n2_adj_140(n2_adj_663), .\read_value[29]_adj_141 (read_value[29]), 
            .n1_adj_142(n1_adj_519), .\read_value[22]_adj_143 (read_value_adj_693[22]), 
            .\read_size[2]_adj_144 (read_size_adj_694[2]), .\read_size[2]_adj_145 (read_size_adj_746[2]), 
            .\read_size[2]_adj_146 (read_size_adj_706[2]), .\read_size[2]_adj_147 (read_size_adj_786[2]), 
            .n4_adj_148(n4_adj_604), .\read_value[3]_adj_149 (read_value_adj_785[3]), 
            .\read_value[3]_adj_150 (read_value_adj_745[3]), .\read_value[3]_adj_151 (read_value[3]), 
            .n2_adj_152(n2_adj_600), .\read_value[31]_adj_153 (read_value[31]), 
            .n1_adj_154(n1_adj_601), .\read_value[31]_adj_155 (read_value_adj_693[31]), 
            .n2_adj_156(n2_adj_442), .n4_adj_157(n4_adj_603), .\read_value[2]_adj_158 (read_value_adj_785[2]), 
            .\read_value[2]_adj_159 (read_value_adj_745[2]), .\read_value[2]_adj_160 (read_value[2]), 
            .\read_value[28]_adj_161 (read_value[28]), .n1_adj_162(n1_adj_649), 
            .\read_value[28]_adj_163 (read_value_adj_693[28]), .n1_adj_164(n1_adj_605), 
            .\read_value[1]_adj_165 (read_value_adj_693[1]), .n6_adj_166(n6_adj_606), 
            .\read_value[1]_adj_167 (read_value_adj_745[1]), .n4_adj_168(n4_adj_602), 
            .\read_value[0]_adj_169 (read_value_adj_785[0]), .\read_value[0]_adj_170 (read_value_adj_745[0]), 
            .\read_value[0]_adj_171 (read_value[0]), .\read_value[29]_adj_172 (read_value_adj_693[29]), 
            .n2_adj_173(n2_adj_591), .n2_adj_174(n2), .\read_value[27]_adj_175 (read_value[27]), 
            .n1_adj_176(n1), .\read_value[21]_adj_177 (read_value[21]), 
            .n1_adj_178(n1_adj_643), .\read_value[27]_adj_179 (read_value_adj_693[27]), 
            .n2_adj_180(n2_adj_394), .\read_value[26]_adj_181 (read_value[26]), 
            .n1_adj_182(n1_adj_395), .\read_value[26]_adj_183 (read_value_adj_693[26]), 
            .\read_value[21]_adj_184 (read_value_adj_693[21]), .n31057(n31057), 
            .debug_c_c(debug_c_c), .n28352(n28352), .GND_net(GND_net), 
            .n32375(n32375), .rc_ch8_c(rc_ch8_c), .n12030(n12030), .n30942(n30942), 
            .n28337(n28337), .n31041(n31041), .rc_ch7_c(rc_ch7_c), .n12031(n12031), 
            .n31025(n31025), .n11987(n11987), .n34347(n34347), .n31050(n31050), 
            .rc_ch4_c(rc_ch4_c), .n30958(n30958), .n28331(n28331), .n12138(n12138), 
            .n28345(n28345), .n30999(n30999), .rc_ch3_c(rc_ch3_c), .n31033(n31033), 
            .n32369(n32369), .n14446(n14446), .n1000(n1000), .n988(n988), 
            .rc_ch2_c(rc_ch2_c), .n54(n54), .n4_adj_185(n4_adj_595), .n32374(n32374), 
            .n31079(n31079), .n28339(n28339), .rc_ch1_c(rc_ch1_c), .n30940(n30940)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(622[15] 634[41])
    \ProtocolInterface(baud_div=12)  protocol_interface (.n32378(n32378), 
            .n30431(n30431), .databus({databus}), .n224({n224}), .n3451({n3451}), 
            .debug_c_c(debug_c_c), .register_addr({register_addr}), .n30418(n30418), 
            .n32420(n32420), .n3363(n3363), .n1318(n1286[0]), .n9(n9_adj_667), 
            .n1304(n1286[14]), .n1310(n1286[8]), .n12098(n12098), .databus_out({databus_out}), 
            .\sendcount[1] (sendcount[1]), .\select[1] (select[1]), .n12788(n12788), 
            .n32472(n32472), .n32395(n32395), .n224_adj_42({n224_adj_789}), 
            .n3181({n3181}), .\select[2] (select[2]), .\select[4] (select[4]), 
            .\select[7] (select[7]), .rw(rw), .\steps_reg[7] (steps_reg[7]), 
            .n9_adj_33(n9), .n4(n4_adj_479), .debug_c_7(debug_c_7), .n32536(n32536), 
            .n11271(n11271), .n5(n5), .n6(n6_adj_592), .\reg_size[2] (reg_size[2]), 
            .n32511(n32511), .n34347(n34347), .n32525(n32525), .n30594(n30594), 
            .n11753(n11753), .\steps_reg[5] (steps_reg_adj_704[5]), .n14(n14_adj_647), 
            .\steps_reg[3] (steps_reg_adj_704[3]), .n15(n15), .\steps_reg[5]_adj_34 (steps_reg_adj_744[5]), 
            .n14_adj_35(n14_adj_598), .\steps_reg[3]_adj_36 (steps_reg_adj_744[3]), 
            .n15_adj_37(n15_adj_440), .\steps_reg[5]_adj_38 (steps_reg_adj_784[5]), 
            .n14_adj_39(n14_adj_662), .\steps_reg[3]_adj_40 (steps_reg_adj_784[3]), 
            .n15_adj_41(n15_adj_659), .debug_c_2(debug_c_2), .debug_c_3(debug_c_3), 
            .debug_c_4(debug_c_4), .debug_c_5(debug_c_5), .n34344(n34344), 
            .\reset_count[14] (reset_count[14]), .\reset_count[12] (reset_count[12]), 
            .\reset_count[13] (reset_count[13]), .n30429(n30429), .\reset_count[10] (reset_count[10]), 
            .\reset_count[9] (reset_count[9]), .n19896(n19896), .n9395(n9395), 
            .GND_net(GND_net), .state({state_adj_832}), .\rdata[0] (rdata[0]), 
            .n29195(n29195), .\rdata[1] (rdata[1]), .n183(n183), .n32(n32), 
            .bclk(bclk), .n31583(n31583), .n32436(n32436), .n32543(n32543), 
            .n32542(n32542), .n32461(n32461), .n9396_c(n9396_c), .n31642(n31642)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[26] 485[57])
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.GND_net(GND_net), .n224({n224}), 
            .n32486(n32486), .n34347(n34347), .n32387(n32387), .n32473(n32473), 
            .n32405(n32405), .rw(rw), .n30450(n30450), .n32420(n32420), 
            .n30283(n30283), .n12434(n12434), .\register_addr[0] (register_addr[0]), 
            .debug_c_c(debug_c_c), .n34351(n34351), .n3451({n3451}), .n34348(n34348), 
            .\read_size[0] (read_size_adj_694[0]), .n11966(n11966), .n30743(n30743), 
            .n34349(n34349), .Stepper_X_M0_c_0(Stepper_X_M0_c_0), .n579(n571[0]), 
            .prev_select(prev_select), .n32435(n32435), .n34350(n34350), 
            .\register_addr[5] (register_addr[5]), .n34344(n34344), .n32378(n32378), 
            .\steps_reg[7] (steps_reg[7]), .n30364(n30364), .limit_c_0(limit_c_0), 
            .n32509(n32509), .n32508(n32508), .n32488(n32488), .n302(n302), 
            .\register_addr[1] (register_addr[1]), .n32527(n32527), .n32453(n32453), 
            .read_value({read_value_adj_693}), .\databus[31] (databus[31]), 
            .n34352(n34352), .\databus[30] (databus[30]), .\databus[29] (databus[29]), 
            .\databus[26] (databus[26]), .\databus[13] (databus[13]), .\databus[11] (databus[11]), 
            .\databus[10] (databus[10]), .\databus[9] (databus[9]), .\databus[7] (databus[7]), 
            .\databus[6] (databus[6]), .\databus[5] (databus[5]), .n608(n580[4]), 
            .n610(n580[2]), .\control_reg[7] (control_reg[7]), .Stepper_X_En_c(Stepper_X_En_c), 
            .n34353(n34353), .Stepper_X_Dir_c(Stepper_X_Dir_c), .\databus[3] (databus[3]), 
            .Stepper_X_M2_c_2(Stepper_X_M2_c_2), .Stepper_X_M1_c_1(Stepper_X_M1_c_1), 
            .\databus[1] (databus[1]), .\read_size[2] (read_size_adj_694[2]), 
            .n32463(n32463), .\register_addr[4] (register_addr[4]), .\register_addr[3] (register_addr[3]), 
            .n11753(n11753), .n30431(n30431), .n18(n18), .\register_addr[6] (register_addr[6]), 
            .\register_addr[7] (register_addr[7]), .n32478(n32478), .\databus[8] (databus[8]), 
            .\databus[12] (databus[12]), .\databus[14] (databus[14]), .\databus[15] (databus[15]), 
            .\databus[16] (databus[16]), .\databus[17] (databus[17]), .\databus[18] (databus[18]), 
            .\databus[19] (databus[19]), .\databus[20] (databus[20]), .\databus[21] (databus[21]), 
            .\databus[22] (databus[22]), .\databus[23] (databus[23]), .n32388(n32388), 
            .n32525(n32525), .n20291(n20291), .n28386(n28386), .\databus[24] (databus[24]), 
            .\databus[25] (databus[25]), .\databus[27] (databus[27]), .\databus[28] (databus[28]), 
            .n11645(n11645), .n32413(n32413), .n30594(n30594), .n8048(n8048), 
            .VCC_net(VCC_net), .Stepper_X_nFault_c(Stepper_X_nFault_c), 
            .Stepper_X_Step_c(Stepper_X_Step_c), .n9(n9), .n28360(n28360)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(559[25] 572[45])
    CCU2D reset_count_2172_2173_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27793), .S0(n66_adj_1126[13]), 
          .S1(n66_adj_1126[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27792), .COUT(n27793), .S0(n66_adj_1126[11]), 
          .S1(n66_adj_1126[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27791), .COUT(n27792), .S0(n66_adj_1126[9]), 
          .S1(n66_adj_1126[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27790), .COUT(n27791), .S0(n66_adj_1126[7]), 
          .S1(n66_adj_1126[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27789), .COUT(n27790), .S0(n66_adj_1126[5]), 
          .S1(n66_adj_1126[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_7.INJECT1_1 = "NO";
    LUT4 Select_3601_i1_2_lut_3_lut_4_lut (.A(n32469), .B(n30454), .C(read_value_adj_785[16]), 
         .D(rw), .Z(n1_adj_641)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3601_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D reset_count_2172_2173_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27788), .COUT(n27789), .S0(n66_adj_1126[3]), 
          .S1(n66_adj_1126[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_5.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27787), .COUT(n27788), .S0(n66_adj_1126[1]), 
          .S1(n66_adj_1126[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27787), .S1(n66_adj_1126[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2172_2173_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2172_2173_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_1.INJECT1_1 = "NO";
    ClockDivider_U10 pwm_clk_div (.debug_c_c(debug_c_c), .n241(n241), .n34347(n34347), 
            .n6674(n6674), .n32375(n32375), .n31079(n31079), .n32374(n32374), 
            .n30942(n30942), .n12030(n12030), .n31025(n31025), .n12031(n12031), 
            .n30958(n30958), .n28331(n28331), .n30940(n30940), .n28339(n28339), 
            .n31033(n31033), .n28345(n28345), .n31041(n31041), .n28337(n28337), 
            .n31057(n31057), .n28352(n28352), .n988(n988), .n6(n6_adj_439), 
            .n30999(n30999), .n12138(n12138), .n31050(n31050), .n11987(n11987), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(508[15] 511[41])
    
endmodule
//
// Verilog Description of module PWMPeripheral
//

module PWMPeripheral (n32478, n32488, rw, n34347, \read_size[0] , 
            debug_c_c, n30743, n34349, \databus[0] , \select[2] , 
            read_value, n282, n34353, \databus[6] , \databus[5] , 
            \databus[4] , \databus[3] , \databus[2] , \databus[1] , 
            n32471, \register_addr[0] , n34344, n64, \count[0] , n32375, 
            motor_pwm_r_c, GND_net, n9633, n14322, \count[1] , \count[2] , 
            \count[3] , \count[4] , \count[5] , \count[6] , \count[7] , 
            \count[8] , n3589, n7893, n7902, n10513, n14473, \count[0]_adj_194 , 
            \count[12] , \count[11] , \count[9] , \count[8]_adj_195 , 
            \count[6]_adj_196 , \count[5]_adj_197 , \count[3]_adj_198 , 
            \count[2]_adj_199 , \count[1]_adj_200 , motor_pwm_l_c, n28488, 
            n32385, n10, n12, \reset_count[6] , n30518, \reset_count[4] , 
            \reset_count[5] , n30519, n3586, n6, \reset_count[8] , 
            \reset_count[7] , n32430, n6_adj_201, n8, n7912, n7906, 
            n7905, n7908, n7910, n7909, n7911) /* synthesis syn_module_defined=1 */ ;
    input n32478;
    input n32488;
    input rw;
    input n34347;
    output \read_size[0] ;
    input debug_c_c;
    input n30743;
    input n34349;
    input \databus[0] ;
    input \select[2] ;
    output [7:0]read_value;
    input n282;
    input n34353;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    input n32471;
    input \register_addr[0] ;
    input n34344;
    output n64;
    output \count[0] ;
    input n32375;
    output motor_pwm_r_c;
    input GND_net;
    output n9633;
    input n14322;
    output \count[1] ;
    output \count[2] ;
    output \count[3] ;
    output \count[4] ;
    output \count[5] ;
    output \count[6] ;
    output \count[7] ;
    output \count[8] ;
    input n3589;
    output [7:0]n7893;
    output n7902;
    output n10513;
    input n14473;
    output \count[0]_adj_194 ;
    output \count[12] ;
    output \count[11] ;
    output \count[9] ;
    output \count[8]_adj_195 ;
    output \count[6]_adj_196 ;
    output \count[5]_adj_197 ;
    output \count[3]_adj_198 ;
    output \count[2]_adj_199 ;
    output \count[1]_adj_200 ;
    output motor_pwm_l_c;
    input n28488;
    output n32385;
    input n10;
    output n12;
    input \reset_count[6] ;
    output n30518;
    input \reset_count[4] ;
    input \reset_count[5] ;
    output n30519;
    input n3586;
    output n6;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n32430;
    input n6_adj_201;
    output n8;
    output n7912;
    output n7906;
    output n7905;
    output n7908;
    output n7910;
    output n7909;
    output n7911;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n32537, n32451, n8052, n12099;
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(55[12:20])
    
    wire n32423, prev_select;
    wire [7:0]n4894;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(55[12:20])
    
    wire n12566, n32424, n20512;
    
    LUT4 i2_3_lut_rep_326_4_lut (.A(n32478), .B(n32488), .C(n32537), .D(rw), 
         .Z(n32451)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_3_lut_rep_326_4_lut.init = 16'h0010;
    LUT4 i2_3_lut_3_lut_4_lut (.A(n32478), .B(n32488), .C(n32537), .D(n34347), 
         .Z(n8052)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i2_3_lut_3_lut_4_lut.init = 16'h00e0;
    FD1P3AX read_size__i1 (.D(n30743), .SP(n12099), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n32423), .PD(n34349), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam prev_select_138.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n4894[1]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n4894[2]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n4894[3]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n4894[4]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n4894[5]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX register_0__i16 (.D(n282), .SP(n12566), .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n32424), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n32424), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n32424), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n32424), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n32424), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n32424), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n32424), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n282), .SP(n20512), .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n32423), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n32423), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n32423), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n32423), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n32423), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n32423), .PD(n34353), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i2.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n4894[6]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n4894[7]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 i24738_2_lut_rep_298_4_lut (.A(rw), .B(n32537), .C(n32471), .D(\register_addr[0] ), 
         .Z(n32423)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i24738_2_lut_rep_298_4_lut.init = 16'h0004;
    LUT4 i3870_2_lut_rep_299_4_lut (.A(rw), .B(n32537), .C(n32471), .D(\register_addr[0] ), 
         .Z(n32424)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3870_2_lut_rep_299_4_lut.init = 16'h0400;
    LUT4 mux_1586_Mux_1_i1_3_lut (.A(\register[0] [1]), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n4894[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_2_i1_3_lut (.A(\register[0] [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n4894[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_3_i1_3_lut (.A(\register[0] [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n4894[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_4_i1_3_lut (.A(\register[0] [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n4894[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_5_i1_3_lut (.A(\register[0] [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n4894[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n4894[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n4894[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_412 (.A(\select[2] ), .B(prev_select), .Z(n32537)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(82[8:29])
    defparam i1_2_lut_rep_412.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\select[2] ), .B(prev_select), .C(n34347), 
         .Z(n12099)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(82[8:29])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 i24731_2_lut_3_lut (.A(\register_addr[0] ), .B(n32451), .C(n34347), 
         .Z(n20512)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(103[9] 108[16])
    defparam i24731_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n32451), .C(n34347), 
         .Z(n12566)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(103[9] 108[16])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    FD1P3IX read_value__i0 (.D(n4894[0]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_1586_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n4894[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 i16_2_lut (.A(\select[2] ), .B(n34344), .Z(n64)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(68[19:32])
    defparam i16_2_lut.init = 16'h8888;
    PWMGenerator right (.count({Open_32, Open_33, Open_34, Open_35, 
            \count[8] , \count[7] , \count[6] , \count[5] , \count[4] , 
            \count[3] , \count[2] , \count[1] , \count[0] }), .debug_c_c(debug_c_c), 
            .n32375(n32375), .motor_pwm_r_c(motor_pwm_r_c), .GND_net(GND_net), 
            .n9633(n9633), .n14322(n14322), .\register[1] ({\register[1] }), 
            .n34347(n34347), .n3589(n3589), .n7893({n7893}), .n7902(n7902)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(118[15] 121[34])
    PWMGenerator_U6 left (.debug_c_c(debug_c_c), .n10513(n10513), .n14473(n14473), 
            .\register[0] ({\register[0] }), .count({\count[12] , \count[11] , 
            Open_36, Open_37, Open_38, Open_39, Open_40, Open_41, 
            Open_42, Open_43, Open_44, Open_45, \count[0]_adj_194 }), 
            .n32375(n32375), .\count[9] (\count[9] ), .\count[8] (\count[8]_adj_195 ), 
            .\count[6] (\count[6]_adj_196 ), .\count[5] (\count[5]_adj_197 ), 
            .\count[3] (\count[3]_adj_198 ), .\count[2] (\count[2]_adj_199 ), 
            .\count[1] (\count[1]_adj_200 ), .n34347(n34347), .motor_pwm_l_c(motor_pwm_l_c), 
            .GND_net(GND_net), .n28488(n28488), .n32385(n32385), .n10(n10), 
            .n12(n12), .\reset_count[6] (\reset_count[6] ), .n30518(n30518), 
            .\reset_count[4] (\reset_count[4] ), .\reset_count[5] (\reset_count[5] ), 
            .n30519(n30519), .n3586(n3586), .n6(n6), .\reset_count[8] (\reset_count[8] ), 
            .\reset_count[7] (\reset_count[7] ), .n32430(n32430), .n6_adj_193(n6_adj_201), 
            .n8(n8), .n7912(n7912), .n7906(n7906), .n7905(n7905), .n7908(n7908), 
            .n7910(n7910), .n7909(n7909), .n7911(n7911)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(114[15] 117[34])
    
endmodule
//
// Verilog Description of module PWMGenerator
//

module PWMGenerator (count, debug_c_c, n32375, motor_pwm_r_c, GND_net, 
            n9633, n14322, \register[1] , n34347, n3589, n7893, 
            n7902) /* synthesis syn_module_defined=1 */ ;
    output [12:0]count;
    input debug_c_c;
    input n32375;
    output motor_pwm_r_c;
    input GND_net;
    output n9633;
    input n14322;
    input [7:0]\register[1] ;
    input n34347;
    input n3589;
    output [7:0]n7893;
    output n7902;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n8031;
    wire [12:0]n43;
    
    wire n28540;
    wire [7:0]latched_width;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(15[12:25])
    wire [12:0]n28;
    wire [12:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    
    wire n30359, n19891, n17, n16, n30626, n8, n27618, n27617, 
        n27616, n27615, n7, n30694, n30757, n30666, n27939, n27938, 
        n27937, n27936, n27935, n27934;
    
    FD1P3IX count__i0 (.D(n43[0]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i0.GSR = "ENABLED";
    OFS1P3DX pwm_19 (.D(n28540), .SP(n32375), .SCLK(debug_c_c), .CD(GND_net), 
            .Q(motor_pwm_r_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam pwm_19.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i0 (.D(\register[1] [0]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i0.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i1 (.D(\register[1] [1]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i1.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n28[1]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n28[2]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n28[3]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n28[4]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n28[5]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n28[6]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n28[7]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n28[8]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n28[9]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n28[10]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i2 (.D(\register[1] [2]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i2.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i3 (.D(\register[1] [3]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i3.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i4 (.D(\register[1] [4]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i4.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i5 (.D(\register[1] [5]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i5.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i6 (.D(\register[1] [6]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i6.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n28[11]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n28[12]), .SP(n32375), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i12.GSR = "ENABLED";
    LUT4 i2274_4_lut (.A(n32375), .B(n30359), .C(n34347), .D(n19891), 
         .Z(n8031)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i2274_4_lut.init = 16'ha0a8;
    LUT4 i9_4_lut (.A(n17), .B(count[5]), .C(n16), .D(n30626), .Z(n30359)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i9_4_lut.init = 16'h0080;
    LUT4 i7_4_lut (.A(count[0]), .B(count_c[9]), .C(count_c[12]), .D(count[6]), 
         .Z(n17)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(count[7]), .B(count[8]), .C(count[3]), .D(count[1]), 
         .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i24272_2_lut (.A(count_c[10]), .B(count_c[11]), .Z(n30626)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24272_2_lut.init = 16'heeee;
    LUT4 i14162_2_lut (.A(count[4]), .B(count[2]), .Z(n19891)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14162_2_lut.init = 16'heeee;
    LUT4 i24773_4_lut (.A(count_c[11]), .B(n3589), .C(count_c[12]), .D(n8), 
         .Z(n28540)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24773_4_lut.init = 16'h0001;
    LUT4 i2_2_lut (.A(count_c[9]), .B(count_c[10]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(26[9:19])
    defparam i2_2_lut.init = 16'heeee;
    FD1P3IX latched_width_i0_i7 (.D(\register[1] [7]), .SP(n9633), .CD(n14322), 
            .CK(debug_c_c), .Q(latched_width[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i7.GSR = "ENABLED";
    CCU2D add_2161_9 (.A0(latched_width[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27618), .S0(n7893[7]), .S1(n7902));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_9.INIT0 = 16'h5555;
    defparam add_2161_9.INIT1 = 16'h0000;
    defparam add_2161_9.INJECT1_0 = "NO";
    defparam add_2161_9.INJECT1_1 = "NO";
    CCU2D add_2161_7 (.A0(latched_width[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27617), .COUT(n27618), .S0(n7893[5]), 
          .S1(n7893[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_7.INIT0 = 16'h5555;
    defparam add_2161_7.INIT1 = 16'h5555;
    defparam add_2161_7.INJECT1_0 = "NO";
    defparam add_2161_7.INJECT1_1 = "NO";
    CCU2D add_2161_5 (.A0(latched_width[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27616), .COUT(n27617), .S0(n7893[3]), 
          .S1(n7893[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_5.INIT0 = 16'h5555;
    defparam add_2161_5.INIT1 = 16'h5555;
    defparam add_2161_5.INJECT1_0 = "NO";
    defparam add_2161_5.INJECT1_1 = "NO";
    CCU2D add_2161_3 (.A0(latched_width[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27615), .COUT(n27616), .S0(n7893[1]), 
          .S1(n7893[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_3.INIT0 = 16'h5555;
    defparam add_2161_3.INIT1 = 16'h5555;
    defparam add_2161_3.INJECT1_0 = "NO";
    defparam add_2161_3.INJECT1_1 = "NO";
    CCU2D add_2161_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(latched_width[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27615), .S1(n7893[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_1.INIT0 = 16'hF000;
    defparam add_2161_1.INIT1 = 16'h5555;
    defparam add_2161_1.INJECT1_0 = "NO";
    defparam add_2161_1.INJECT1_1 = "NO";
    LUT4 i4_4_lut (.A(n7), .B(n30626), .C(n19891), .D(count[0]), .Z(n9633)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h0002;
    LUT4 i2_4_lut (.A(n30694), .B(n32375), .C(n30757), .D(n30666), .Z(n7)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0004;
    LUT4 i24337_2_lut (.A(count_c[9]), .B(count[3]), .Z(n30694)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24337_2_lut.init = 16'heeee;
    LUT4 i24399_4_lut (.A(count[7]), .B(count[5]), .C(count[1]), .D(count_c[12]), 
         .Z(n30757)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24399_4_lut.init = 16'hfffe;
    LUT4 i24312_2_lut (.A(count[6]), .B(count[8]), .Z(n30666)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24312_2_lut.init = 16'heeee;
    CCU2D add_9_13 (.A0(count_c[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27939), .S0(n28[11]), .S1(n28[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_13.INIT0 = 16'h5aaa;
    defparam add_9_13.INIT1 = 16'h5aaa;
    defparam add_9_13.INJECT1_0 = "NO";
    defparam add_9_13.INJECT1_1 = "NO";
    CCU2D add_9_11 (.A0(count_c[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27938), .COUT(n27939), .S0(n28[9]), .S1(n28[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_11.INIT0 = 16'h5aaa;
    defparam add_9_11.INIT1 = 16'h5aaa;
    defparam add_9_11.INJECT1_0 = "NO";
    defparam add_9_11.INJECT1_1 = "NO";
    CCU2D add_9_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27937), 
          .COUT(n27938), .S0(n28[7]), .S1(n28[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_9.INIT0 = 16'h5aaa;
    defparam add_9_9.INIT1 = 16'h5aaa;
    defparam add_9_9.INJECT1_0 = "NO";
    defparam add_9_9.INJECT1_1 = "NO";
    CCU2D add_9_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27936), 
          .COUT(n27937), .S0(n28[5]), .S1(n28[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_7.INIT0 = 16'h5aaa;
    defparam add_9_7.INIT1 = 16'h5aaa;
    defparam add_9_7.INJECT1_0 = "NO";
    defparam add_9_7.INJECT1_1 = "NO";
    CCU2D add_9_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27935), 
          .COUT(n27936), .S0(n28[3]), .S1(n28[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_5.INIT0 = 16'h5aaa;
    defparam add_9_5.INIT1 = 16'h5aaa;
    defparam add_9_5.INJECT1_0 = "NO";
    defparam add_9_5.INJECT1_1 = "NO";
    CCU2D add_9_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27934), 
          .COUT(n27935), .S0(n28[1]), .S1(n28[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_3.INIT0 = 16'h5aaa;
    defparam add_9_3.INIT1 = 16'h5aaa;
    defparam add_9_3.INJECT1_0 = "NO";
    defparam add_9_3.INJECT1_1 = "NO";
    CCU2D add_9_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27934), 
          .S1(n43[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_1.INIT0 = 16'hF000;
    defparam add_9_1.INIT1 = 16'h5555;
    defparam add_9_1.INJECT1_0 = "NO";
    defparam add_9_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMGenerator_U6
//

module PWMGenerator_U6 (debug_c_c, n10513, n14473, \register[0] , count, 
            n32375, \count[9] , \count[8] , \count[6] , \count[5] , 
            \count[3] , \count[2] , \count[1] , n34347, motor_pwm_l_c, 
            GND_net, n28488, n32385, n10, n12, \reset_count[6] , 
            n30518, \reset_count[4] , \reset_count[5] , n30519, n3586, 
            n6, \reset_count[8] , \reset_count[7] , n32430, n6_adj_193, 
            n8, n7912, n7906, n7905, n7908, n7910, n7909, n7911) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output n10513;
    input n14473;
    input [7:0]\register[0] ;
    output [12:0]count;
    input n32375;
    output \count[9] ;
    output \count[8] ;
    output \count[6] ;
    output \count[5] ;
    output \count[3] ;
    output \count[2] ;
    output \count[1] ;
    input n34347;
    output motor_pwm_l_c;
    input GND_net;
    input n28488;
    output n32385;
    input n10;
    output n12;
    input \reset_count[6] ;
    output n30518;
    input \reset_count[4] ;
    input \reset_count[5] ;
    output n30519;
    input n3586;
    output n6;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n32430;
    input n6_adj_193;
    output n8;
    output n7912;
    output n7906;
    output n7905;
    output n7908;
    output n7910;
    output n7909;
    output n7911;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [7:0]latched_width;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(15[12:25])
    wire [12:0]n42;
    
    wire n8027;
    wire [12:0]n43;
    wire [12:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    wire [12:0]n28;
    
    wire n28566, n30620, n15_adj_382, n14;
    wire [7:0]n7903;
    
    wire n32512, n30747, n30783, n30749, n27932, n27931, n27930, 
        n27929, n27928, n27927, n27926, n27925, n27924, n27923;
    
    FD1P3JX latched_width_i0_i2 (.D(\register[0] [2]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i2.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i1 (.D(\register[0] [1]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i1.GSR = "ENABLED";
    FD1P3AX count__i0 (.D(n42[0]), .SP(n32375), .CK(debug_c_c), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n43[12]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n43[11]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n43[10]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(count_c[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n43[9]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n43[8]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n43[7]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(count_c[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n43[6]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n43[5]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n43[4]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(count_c[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n43[3]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[3] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n43[2]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[2] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n43[1]), .SP(n32375), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i14029_2_lut (.A(n28[0]), .B(n8027), .Z(n42[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i14029_2_lut.init = 16'h2222;
    LUT4 i2270_4_lut (.A(n32375), .B(n28566), .C(n34347), .D(n30620), 
         .Z(n8027)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i2270_4_lut.init = 16'ha0a8;
    LUT4 i8_4_lut (.A(n15_adj_382), .B(\count[8] ), .C(n14), .D(\count[9] ), 
         .Z(n28566)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(\count[5] ), .B(\count[6] ), .C(count[0]), .D(\count[1] ), 
         .Z(n15_adj_382)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(count[12]), .B(count_c[7]), .C(\count[3] ), .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    FD1P3JX latched_width_i0_i0 (.D(\register[0] [0]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i0.GSR = "ENABLED";
    FD1P3IX pwm_19 (.D(n28488), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(motor_pwm_l_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam pwm_19.GSR = "ENABLED";
    LUT4 i10_2_lut_rep_260 (.A(n7903[7]), .B(count_c[7]), .Z(n32385)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam i10_2_lut_rep_260.init = 16'h6666;
    LUT4 LessThan_1434_i12_3_lut_3_lut (.A(n7903[7]), .B(count_c[7]), .C(n10), 
         .Z(n12)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam LessThan_1434_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i45_2_lut_rep_387 (.A(\count[2] ), .B(count_c[4]), .Z(n32512)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i45_2_lut_rep_387.init = 16'heeee;
    LUT4 i24266_3_lut_4_lut (.A(\count[2] ), .B(count_c[4]), .C(count[11]), 
         .D(count_c[10]), .Z(n30620)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24266_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n32375), .B(n32512), .C(n30747), .D(n30783), .Z(n10513)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0002;
    LUT4 i24389_4_lut (.A(count[11]), .B(count_c[7]), .C(\count[5] ), 
         .D(\count[9] ), .Z(n30747)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24389_4_lut.init = 16'hfffe;
    LUT4 i24425_4_lut (.A(count[12]), .B(n30749), .C(\count[8] ), .D(count[0]), 
         .Z(n30783)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24425_4_lut.init = 16'hfffe;
    LUT4 i24391_4_lut (.A(\count[3] ), .B(count_c[10]), .C(\count[1] ), 
         .D(\count[6] ), .Z(n30749)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24391_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(\reset_count[6] ), .B(n30518), .C(\reset_count[4] ), 
         .D(\reset_count[5] ), .Z(n30519)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'heeec;
    LUT4 i1_2_lut (.A(count_c[10]), .B(n3586), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(26[9:19])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_470 (.A(\reset_count[8] ), .B(\reset_count[7] ), .Z(n30518)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_470.init = 16'heeee;
    FD1P3IX latched_width_i0_i7 (.D(\register[0] [7]), .SP(n10513), .CD(n14473), 
            .CK(debug_c_c), .Q(latched_width[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i7.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i6 (.D(\register[0] [6]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i6.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i5 (.D(\register[0] [5]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i5.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i4 (.D(\register[0] [4]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i4.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i3 (.D(\register[0] [3]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i3.GSR = "ENABLED";
    LUT4 i9_2_lut_rep_305 (.A(n7903[4]), .B(count_c[4]), .Z(n32430)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam i9_2_lut_rep_305.init = 16'h6666;
    LUT4 LessThan_1434_i8_3_lut_3_lut (.A(n7903[4]), .B(count_c[4]), .C(n6_adj_193), 
         .Z(n8)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam LessThan_1434_i8_3_lut_3_lut.init = 16'hd4d4;
    CCU2D add_9_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27932), .S0(n43[11]), .S1(n43[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_13.INIT0 = 16'h5aaa;
    defparam add_9_13.INIT1 = 16'h5aaa;
    defparam add_9_13.INJECT1_0 = "NO";
    defparam add_9_13.INJECT1_1 = "NO";
    CCU2D add_9_11 (.A0(\count[9] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27931), .COUT(n27932), .S0(n43[9]), .S1(n43[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_11.INIT0 = 16'h5aaa;
    defparam add_9_11.INIT1 = 16'h5aaa;
    defparam add_9_11.INJECT1_0 = "NO";
    defparam add_9_11.INJECT1_1 = "NO";
    CCU2D add_9_9 (.A0(count_c[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27930), .COUT(n27931), .S0(n43[7]), .S1(n43[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_9.INIT0 = 16'h5aaa;
    defparam add_9_9.INIT1 = 16'h5aaa;
    defparam add_9_9.INJECT1_0 = "NO";
    defparam add_9_9.INJECT1_1 = "NO";
    CCU2D add_9_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27929), .COUT(n27930), .S0(n43[5]), .S1(n43[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_7.INIT0 = 16'h5aaa;
    defparam add_9_7.INIT1 = 16'h5aaa;
    defparam add_9_7.INJECT1_0 = "NO";
    defparam add_9_7.INJECT1_1 = "NO";
    CCU2D add_9_5 (.A0(\count[3] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27928), .COUT(n27929), .S0(n43[3]), .S1(n43[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_5.INIT0 = 16'h5aaa;
    defparam add_9_5.INIT1 = 16'h5aaa;
    defparam add_9_5.INJECT1_0 = "NO";
    defparam add_9_5.INJECT1_1 = "NO";
    CCU2D add_9_3 (.A0(\count[1] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[2] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27927), .COUT(n27928), .S0(n43[1]), .S1(n43[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_3.INIT0 = 16'h5aaa;
    defparam add_9_3.INIT1 = 16'h5aaa;
    defparam add_9_3.INJECT1_0 = "NO";
    defparam add_9_3.INJECT1_1 = "NO";
    CCU2D add_9_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27927), 
          .S1(n28[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_1.INIT0 = 16'hF000;
    defparam add_9_1.INIT1 = 16'h5555;
    defparam add_9_1.INJECT1_0 = "NO";
    defparam add_9_1.INJECT1_1 = "NO";
    CCU2D add_2162_9 (.A0(latched_width[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27926), .S0(n7903[7]), .S1(n7912));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_9.INIT0 = 16'h5555;
    defparam add_2162_9.INIT1 = 16'h0000;
    defparam add_2162_9.INJECT1_0 = "NO";
    defparam add_2162_9.INJECT1_1 = "NO";
    CCU2D add_2162_7 (.A0(latched_width[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27925), .COUT(n27926), .S0(n7906), .S1(n7905));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_7.INIT0 = 16'h5555;
    defparam add_2162_7.INIT1 = 16'h5555;
    defparam add_2162_7.INJECT1_0 = "NO";
    defparam add_2162_7.INJECT1_1 = "NO";
    CCU2D add_2162_5 (.A0(latched_width[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27924), .COUT(n27925), .S0(n7908), .S1(n7903[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_5.INIT0 = 16'h5555;
    defparam add_2162_5.INIT1 = 16'h5555;
    defparam add_2162_5.INJECT1_0 = "NO";
    defparam add_2162_5.INJECT1_1 = "NO";
    CCU2D add_2162_3 (.A0(latched_width[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27923), .COUT(n27924), .S0(n7910), .S1(n7909));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_3.INIT0 = 16'h5555;
    defparam add_2162_3.INIT1 = 16'h5555;
    defparam add_2162_3.INJECT1_0 = "NO";
    defparam add_2162_3.INJECT1_1 = "NO";
    CCU2D add_2162_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(latched_width[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27923), .S1(n7911));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_1.INIT0 = 16'hF000;
    defparam add_2162_1.INIT1 = 16'h5555;
    defparam add_2162_1.INJECT1_0 = "NO";
    defparam add_2162_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (read_value, debug_c_c, n32413, register_addr, 
            n32486, n8048, n11753, n30418, read_size, n302, \register[2] , 
            n34348, \select[1] , \select[4] , n32527, n32469, n32454, 
            n34350, n34349, \register[2][3] , n28386, n32453, n32463, 
            n15, n32462, n4, n10513, n14473, signal_light_c, n9633, 
            n14322, \control_reg[7] , n28360, n18, \control_reg[7]_adj_188 , 
            n28299, stepping, \control_reg[7]_adj_189 , n28401, stepping_adj_190, 
            \control_reg[7]_adj_191 , n28214, stepping_adj_192, rw, 
            n32503, n6, n32478, n11645, \databus[1] , n34347, n32525, 
            xbee_pause_c, n20291, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    output n32413;
    input [7:0]register_addr;
    output n32486;
    input n8048;
    input n11753;
    output n30418;
    output [2:0]read_size;
    input n302;
    output [31:0]\register[2] ;
    input n34348;
    input \select[1] ;
    input \select[4] ;
    input n32527;
    output n32469;
    input n32454;
    input n34350;
    input n34349;
    output \register[2][3] ;
    input n28386;
    input n32453;
    input n32463;
    input n15;
    input n32462;
    input n4;
    input n10513;
    output n14473;
    output signal_light_c;
    input n9633;
    output n14322;
    input \control_reg[7] ;
    input n28360;
    output n18;
    input \control_reg[7]_adj_188 ;
    input n28299;
    output stepping;
    input \control_reg[7]_adj_189 ;
    input n28401;
    output stepping_adj_190;
    input \control_reg[7]_adj_191 ;
    input n28214;
    output stepping_adj_192;
    input rw;
    output n32503;
    output n6;
    input n32478;
    input n11645;
    input \databus[1] ;
    input n34347;
    output n32525;
    input xbee_pause_c;
    output n20291;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30445, n29676, n29675, n29682, n29672, n29664, n29659, 
        n29680, n29685, n29658, n29679, n29677, n29684, n29667, 
        n29666, n29660, n29662, n29674, n29673, n29663, n29671, 
        n29668, n29681, n29683, n29661, n29670, n29678, n29669, 
        n29665, n30444, n32367;
    wire [31:0]read_value_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    
    wire n32368, n7999;
    wire [31:0]n100;
    
    wire prev_clk_1Hz, clk_1Hz;
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n178, prev_select, n27, n16;
    wire [31:0]\register[2]_c ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n32538, force_pause, n21, n14414, n14413, n24, n11, n27_adj_380, 
        n16_adj_381, n28027, n30230, n32510, n27598, n27597, n27596, 
        n27595, n27594, n27593, n27592, n27591, n27590, n27589, 
        n27588, n27587, n27586, n27585, n27584, n27583;
    
    FD1P3AX read_value__i0 (.D(n30445), .SP(n32413), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_361_3_lut_4_lut (.A(register_addr[7]), .B(register_addr[6]), 
         .C(register_addr[5]), .D(register_addr[4]), .Z(n32486)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_361_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX read_value__i31 (.D(n29676), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n29675), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n29682), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n29672), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n29664), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n29659), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n29680), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n29685), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n29658), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n29679), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n29677), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n29684), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n29667), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n29666), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n29660), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n29662), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i16.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(n11753), .B(register_addr[3]), .Z(n30418)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam i1_2_lut.init = 16'h2222;
    FD1P3IX read_value__i15 (.D(n29674), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n29673), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n29663), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n29671), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n29668), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n29681), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n29683), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n29661), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n29670), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n29678), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n29669), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n29665), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n30444), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n32367), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n32368), .SP(n32413), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value_c[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n302), .SP(n32413), .CK(debug_c_c), .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n7999), .CD(n34348), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_149 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_clk_1Hz_149.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_150 (.D(n178), .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam xbee_pause_latched_150.GSR = "ENABLED";
    FD1S3AX prev_select_148 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_select_148.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(register_addr[7]), .B(register_addr[6]), 
         .C(\select[4] ), .D(n32527), .Z(n32469)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'h0010;
    LUT4 n27_bdd_4_lut (.A(n27), .B(n16), .C(register_addr[1]), .D(n32454), 
         .Z(n32368)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n27_bdd_4_lut.init = 16'h00ca;
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n7999), .CD(n34350), 
            .CK(debug_c_c), .Q(\register[2]_c [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n7999), .CD(n34348), 
            .CK(debug_c_c), .Q(\register[2]_c [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n7999), .CD(n34348), 
            .CK(debug_c_c), .Q(\register[2]_c [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n7999), .CD(n34348), 
            .CK(debug_c_c), .Q(\register[2]_c [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n7999), .CD(n34348), 
            .CK(debug_c_c), .Q(\register[2]_c [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n32538), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n7999), .CD(n34349), 
            .CK(debug_c_c), .Q(\register[2]_c [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n7999), .CD(n34348), 
            .CK(debug_c_c), .Q(\register[2]_c [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n7999), .CD(n34349), .CK(debug_c_c), 
            .Q(\register[2]_c [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n7999), .CD(n34348), .CK(debug_c_c), 
            .Q(\register[2]_c [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n7999), .CD(n34349), .CK(debug_c_c), 
            .Q(\register[2]_c [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n7999), .CD(n34349), .CK(debug_c_c), 
            .Q(\register[2]_c [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n7999), .CD(n34349), .CK(debug_c_c), 
            .Q(\register[2]_c [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n7999), .CD(n34349), .CK(debug_c_c), 
            .Q(\register[2]_c [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n7999), .CD(n34348), .CK(debug_c_c), 
            .Q(\register[2][3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(register_addr[2]), 
         .D(register_addr[3]), .Z(n21)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h00fe;
    FD1P3IX read_size_i0_i1 (.D(n28386), .SP(n32413), .CD(n14414), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n32453), .SP(n32413), .CD(n14413), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n7999), .CD(n32463), .CK(debug_c_c), 
            .Q(\register[2]_c [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n7999), .CD(n32463), .CK(debug_c_c), 
            .Q(\register[2]_c [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    PFUMX i33 (.BLUT(n21), .ALUT(n15), .C0(register_addr[1]), .Z(n24));
    LUT4 i1_4_lut (.A(n11), .B(n32462), .C(n4), .D(register_addr[1]), 
         .Z(n30444)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h3022;
    LUT4 i1_2_lut_adj_433 (.A(register_addr[3]), .B(register_addr[2]), .Z(n11)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam i1_2_lut_adj_433.init = 16'h4444;
    LUT4 i8712_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(n10513), 
         .Z(n14473)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i8712_2_lut_3_lut.init = 16'he0e0;
    LUT4 i13950_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(clk_1Hz), 
         .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i13950_2_lut_3_lut.init = 16'hfefe;
    LUT4 i8679_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(n9633), 
         .Z(n14322)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i8679_2_lut_3_lut.init = 16'he0e0;
    LUT4 i2_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(\control_reg[7] ), 
         .D(n28360), .Z(n18)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_434 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_188 ), .D(n28299), .Z(stepping)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_434.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_435 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_189 ), .D(n28401), .Z(stepping_adj_190)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_435.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_436 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_191 ), .D(n28214), .Z(stepping_adj_192)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_436.init = 16'h1000;
    LUT4 i14_2_lut_rep_378 (.A(\select[1] ), .B(rw), .Z(n32503)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam i14_2_lut_rep_378.init = 16'h8888;
    LUT4 Select_3624_i6_2_lut_3_lut (.A(\select[1] ), .B(rw), .C(read_value_c[1]), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam Select_3624_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 n27_bdd_4_lut_adj_437 (.A(n27_adj_380), .B(n16_adj_381), .C(register_addr[1]), 
         .D(n32454), .Z(n32367)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n27_bdd_4_lut_adj_437.init = 16'h00ca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32478), .B(n32527), .C(\register[2]_c [6]), 
         .D(n11645), .Z(n29678)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_438 (.A(n32478), .B(n32527), .C(\register[2]_c [31]), 
         .D(n11645), .Z(n29676)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_438.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_439 (.A(n32478), .B(n32527), .C(\register[2]_c [4]), 
         .D(n11645), .Z(n29665)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_439.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_440 (.A(n32478), .B(n32527), .C(\register[2]_c [8]), 
         .D(n11645), .Z(n29661)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_440.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_441 (.A(n32478), .B(n32527), .C(\register[2]_c [9]), 
         .D(n11645), .Z(n29683)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_441.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_442 (.A(n32478), .B(n32527), .C(\register[2]_c [10]), 
         .D(n11645), .Z(n29681)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_442.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_443 (.A(n32478), .B(n32527), .C(\register[2]_c [11]), 
         .D(n11645), .Z(n29668)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_443.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_444 (.A(n32478), .B(n32527), .C(\register[2]_c [12]), 
         .D(n11645), .Z(n29671)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_444.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_445 (.A(n32478), .B(n32527), .C(\register[2]_c [13]), 
         .D(n11645), .Z(n29663)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_445.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_446 (.A(n32478), .B(n32527), .C(\register[2]_c [14]), 
         .D(n11645), .Z(n29673)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_446.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_447 (.A(n32478), .B(n32527), .C(\register[2]_c [15]), 
         .D(n11645), .Z(n29674)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_447.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_448 (.A(n32478), .B(n32527), .C(\register[2]_c [17]), 
         .D(n11645), .Z(n29660)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_448.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_449 (.A(n32478), .B(n32527), .C(\register[2]_c [18]), 
         .D(n11645), .Z(n29666)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_449.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_450 (.A(n32478), .B(n32527), .C(\register[2]_c [19]), 
         .D(n11645), .Z(n29667)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_450.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_451 (.A(n32478), .B(n32527), .C(\register[2]_c [20]), 
         .D(n11645), .Z(n29684)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_451.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_452 (.A(n32478), .B(n32527), .C(\register[2]_c [30]), 
         .D(n11645), .Z(n29675)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_452.init = 16'h1000;
    FD1P3IX force_pause_151 (.D(\databus[1] ), .SP(n28027), .CD(n32463), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam force_pause_151.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_453 (.A(n32478), .B(n32527), .C(\register[2]_c [21]), 
         .D(n11645), .Z(n29677)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_453.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_454 (.A(n32478), .B(n32527), .C(\register[2]_c [22]), 
         .D(n11645), .Z(n29679)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_454.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_455 (.A(n32478), .B(n32527), .C(\register[2]_c [23]), 
         .D(n11645), .Z(n29658)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_455.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_456 (.A(n32478), .B(n32527), .C(\register[2]_c [24]), 
         .D(n11645), .Z(n29685)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_456.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_457 (.A(n32478), .B(n32527), .C(\register[2]_c [25]), 
         .D(n11645), .Z(n29680)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_457.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_458 (.A(n32478), .B(n32527), .C(\register[2]_c [26]), 
         .D(n11645), .Z(n29659)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_458.init = 16'h1000;
    LUT4 i1_3_lut_4_lut (.A(n32478), .B(n32527), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n30230)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1101;
    LUT4 i1_2_lut_3_lut_4_lut_adj_459 (.A(n32478), .B(n32527), .C(\register[2]_c [29]), 
         .D(n11645), .Z(n29682)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_459.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_460 (.A(n32478), .B(n32527), .C(\register[2]_c [27]), 
         .D(n11645), .Z(n29664)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_460.init = 16'h1000;
    LUT4 i117_2_lut_rep_385 (.A(prev_select), .B(\select[1] ), .Z(n32510)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i117_2_lut_rep_385.init = 16'h4444;
    LUT4 i8648_2_lut_3_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(n30230), .D(n34347), .Z(n14414)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i8648_2_lut_3_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i8647_2_lut_3_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(n30230), .D(n34347), .Z(n14413)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i8647_2_lut_3_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i889_2_lut_rep_288_2_lut_3_lut (.A(prev_select), .B(\select[1] ), 
         .C(n34347), .Z(n32413)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i889_2_lut_rep_288_2_lut_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_3_lut_4_lut_adj_461 (.A(n32478), .B(n32527), .C(\register[2]_c [5]), 
         .D(n11645), .Z(n29669)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_461.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_462 (.A(n32478), .B(n32527), .C(\register[2]_c [7]), 
         .D(n11645), .Z(n29670)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_462.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_463 (.A(n32478), .B(n32527), .C(\register[2]_c [16]), 
         .D(n11645), .Z(n29662)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_463.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_464 (.A(n32478), .B(n32527), .C(\register[2]_c [28]), 
         .D(n11645), .Z(n29672)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_464.init = 16'h1000;
    LUT4 i13835_2_lut_rep_400 (.A(register_addr[7]), .B(register_addr[6]), 
         .Z(n32525)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13835_2_lut_rep_400.init = 16'heeee;
    LUT4 i114_1_lut (.A(xbee_pause_c), .Z(n178)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(54[26:39])
    defparam i114_1_lut.init = 16'h5555;
    LUT4 i14556_3_lut (.A(register_addr[2]), .B(register_addr[1]), .C(register_addr[0]), 
         .Z(n20291)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i14556_3_lut.init = 16'ha8a8;
    LUT4 i1_3_lut_4_lut_adj_465 (.A(register_addr[0]), .B(n32478), .C(n24), 
         .D(n8048), .Z(n30445)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_465.init = 16'h0010;
    LUT4 i1_2_lut_adj_466 (.A(\register[2]_c [2]), .B(register_addr[0]), 
         .Z(n16_adj_381)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_466.init = 16'h2222;
    LUT4 i1_2_lut_adj_467 (.A(\register[2]_c [1]), .B(register_addr[0]), 
         .Z(n16)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_467.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_adj_468 (.A(register_addr[3]), .B(register_addr[2]), 
         .C(\register[0] [2]), .D(register_addr[0]), .Z(n27_adj_380)) /* synthesis lut_function=(A (C+(D))+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_468.init = 16'hffb0;
    LUT4 i1_3_lut_4_lut_adj_469 (.A(register_addr[3]), .B(register_addr[2]), 
         .C(force_pause), .D(register_addr[0]), .Z(n27)) /* synthesis lut_function=(A (C+(D))+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_469.init = 16'hffb0;
    LUT4 i134_2_lut_rep_413 (.A(prev_clk_1Hz), .B(clk_1Hz), .Z(n32538)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i134_2_lut_rep_413.init = 16'h4444;
    LUT4 i2256_2_lut_3_lut (.A(prev_clk_1Hz), .B(clk_1Hz), .C(n34347), 
         .Z(n7999)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i2256_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i2_4_lut (.A(n34347), .B(rw), .C(n32510), .D(n32453), .Z(n28027)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam i2_4_lut.init = 16'h0032;
    CCU2D add_134_33 (.A0(\register[2]_c [31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27598), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_33.INIT0 = 16'h5aaa;
    defparam add_134_33.INIT1 = 16'h0000;
    defparam add_134_33.INJECT1_0 = "NO";
    defparam add_134_33.INJECT1_1 = "NO";
    CCU2D add_134_31 (.A0(\register[2]_c [29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27597), .COUT(n27598), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_31.INIT0 = 16'h5aaa;
    defparam add_134_31.INIT1 = 16'h5aaa;
    defparam add_134_31.INJECT1_0 = "NO";
    defparam add_134_31.INJECT1_1 = "NO";
    CCU2D add_134_29 (.A0(\register[2]_c [27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27596), .COUT(n27597), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_29.INIT0 = 16'h5aaa;
    defparam add_134_29.INIT1 = 16'h5aaa;
    defparam add_134_29.INJECT1_0 = "NO";
    defparam add_134_29.INJECT1_1 = "NO";
    CCU2D add_134_27 (.A0(\register[2]_c [25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27595), .COUT(n27596), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_27.INIT0 = 16'h5aaa;
    defparam add_134_27.INIT1 = 16'h5aaa;
    defparam add_134_27.INJECT1_0 = "NO";
    defparam add_134_27.INJECT1_1 = "NO";
    CCU2D add_134_25 (.A0(\register[2]_c [23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27594), .COUT(n27595), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_25.INIT0 = 16'h5aaa;
    defparam add_134_25.INIT1 = 16'h5aaa;
    defparam add_134_25.INJECT1_0 = "NO";
    defparam add_134_25.INJECT1_1 = "NO";
    CCU2D add_134_23 (.A0(\register[2]_c [21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27593), .COUT(n27594), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_23.INIT0 = 16'h5aaa;
    defparam add_134_23.INIT1 = 16'h5aaa;
    defparam add_134_23.INJECT1_0 = "NO";
    defparam add_134_23.INJECT1_1 = "NO";
    CCU2D add_134_21 (.A0(\register[2]_c [19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27592), .COUT(n27593), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_21.INIT0 = 16'h5aaa;
    defparam add_134_21.INIT1 = 16'h5aaa;
    defparam add_134_21.INJECT1_0 = "NO";
    defparam add_134_21.INJECT1_1 = "NO";
    CCU2D add_134_19 (.A0(\register[2]_c [17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27591), .COUT(n27592), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_19.INIT0 = 16'h5aaa;
    defparam add_134_19.INIT1 = 16'h5aaa;
    defparam add_134_19.INJECT1_0 = "NO";
    defparam add_134_19.INJECT1_1 = "NO";
    CCU2D add_134_17 (.A0(\register[2]_c [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27590), .COUT(n27591), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_17.INIT0 = 16'h5aaa;
    defparam add_134_17.INIT1 = 16'h5aaa;
    defparam add_134_17.INJECT1_0 = "NO";
    defparam add_134_17.INJECT1_1 = "NO";
    CCU2D add_134_15 (.A0(\register[2]_c [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27589), .COUT(n27590), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_15.INIT0 = 16'h5aaa;
    defparam add_134_15.INIT1 = 16'h5aaa;
    defparam add_134_15.INJECT1_0 = "NO";
    defparam add_134_15.INJECT1_1 = "NO";
    CCU2D add_134_13 (.A0(\register[2]_c [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27588), .COUT(n27589), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_13.INIT0 = 16'h5aaa;
    defparam add_134_13.INIT1 = 16'h5aaa;
    defparam add_134_13.INJECT1_0 = "NO";
    defparam add_134_13.INJECT1_1 = "NO";
    CCU2D add_134_11 (.A0(\register[2]_c [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27587), .COUT(n27588), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_11.INIT0 = 16'h5aaa;
    defparam add_134_11.INIT1 = 16'h5aaa;
    defparam add_134_11.INJECT1_0 = "NO";
    defparam add_134_11.INJECT1_1 = "NO";
    CCU2D add_134_9 (.A0(\register[2]_c [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27586), .COUT(n27587), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_9.INIT0 = 16'h5aaa;
    defparam add_134_9.INIT1 = 16'h5aaa;
    defparam add_134_9.INJECT1_0 = "NO";
    defparam add_134_9.INJECT1_1 = "NO";
    CCU2D add_134_7 (.A0(\register[2]_c [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27585), .COUT(n27586), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_7.INIT0 = 16'h5aaa;
    defparam add_134_7.INIT1 = 16'h5aaa;
    defparam add_134_7.INJECT1_0 = "NO";
    defparam add_134_7.INJECT1_1 = "NO";
    CCU2D add_134_5 (.A0(\register[2][3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27584), .COUT(n27585), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_5.INIT0 = 16'h5aaa;
    defparam add_134_5.INIT1 = 16'h5aaa;
    defparam add_134_5.INJECT1_0 = "NO";
    defparam add_134_5.INJECT1_1 = "NO";
    CCU2D add_134_3 (.A0(\register[2]_c [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27583), .COUT(n27584), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_3.INIT0 = 16'h5aaa;
    defparam add_134_3.INIT1 = 16'h5aaa;
    defparam add_134_3.INJECT1_0 = "NO";
    defparam add_134_3.INJECT1_1 = "NO";
    CCU2D add_134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27583), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_1.INIT0 = 16'hF000;
    defparam add_134_1.INIT1 = 16'h5555;
    defparam add_134_1.INJECT1_0 = "NO";
    defparam add_134_1.INJECT1_1 = "NO";
    \ClockDividerP(factor=12000000)  uptime_div (.debug_c_c(debug_c_c), .clk_1Hz(clk_1Hz), 
            .n32463(n32463), .n34347(n34347), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(107[28] 109[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (debug_c_c, clk_1Hz, n32463, n34347, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output clk_1Hz;
    input n32463;
    input n34347;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n2595;
    wire [31:0]n134;
    
    wire n6778, n30948, n27, n28180, n25, n26, n24, n19, n32, 
        n28, n20, n29, n26_adj_374, n27952, n27951, n27950, n27949, 
        n27948, n27947, n27946, n27945, n27944, n27943, n27942, 
        n27941, n27858, n27857, n27856, n27855, n27854, n27853, 
        n27852, n27851, n27850, n27849, n27848, n27847, n27846, 
        n27845, n27844, n27843;
    
    FD1S3IX count_2175__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2595), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i0.GSR = "ENABLED";
    FD1S3IX clk_o_14 (.D(n6778), .CK(debug_c_c), .CD(n32463), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2175__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2595), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i1.GSR = "ENABLED";
    FD1S3IX count_2175__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2595), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i2.GSR = "ENABLED";
    FD1S3IX count_2175__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2595), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i3.GSR = "ENABLED";
    FD1S3IX count_2175__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2595), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i4.GSR = "ENABLED";
    FD1S3IX count_2175__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2595), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i5.GSR = "ENABLED";
    FD1S3IX count_2175__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2595), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i6.GSR = "ENABLED";
    FD1S3IX count_2175__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2595), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i7.GSR = "ENABLED";
    FD1S3IX count_2175__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2595), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i8.GSR = "ENABLED";
    FD1S3IX count_2175__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2595), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i9.GSR = "ENABLED";
    FD1S3IX count_2175__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i10.GSR = "ENABLED";
    FD1S3IX count_2175__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i11.GSR = "ENABLED";
    FD1S3IX count_2175__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i12.GSR = "ENABLED";
    FD1S3IX count_2175__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i13.GSR = "ENABLED";
    FD1S3IX count_2175__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i14.GSR = "ENABLED";
    FD1S3IX count_2175__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i15.GSR = "ENABLED";
    FD1S3IX count_2175__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i16.GSR = "ENABLED";
    FD1S3IX count_2175__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i17.GSR = "ENABLED";
    FD1S3IX count_2175__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i18.GSR = "ENABLED";
    FD1S3IX count_2175__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i19.GSR = "ENABLED";
    FD1S3IX count_2175__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i20.GSR = "ENABLED";
    FD1S3IX count_2175__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i21.GSR = "ENABLED";
    FD1S3IX count_2175__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i22.GSR = "ENABLED";
    FD1S3IX count_2175__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i23.GSR = "ENABLED";
    FD1S3IX count_2175__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i24.GSR = "ENABLED";
    FD1S3IX count_2175__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i25.GSR = "ENABLED";
    FD1S3IX count_2175__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i26.GSR = "ENABLED";
    FD1S3IX count_2175__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i27.GSR = "ENABLED";
    FD1S3IX count_2175__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i28.GSR = "ENABLED";
    FD1S3IX count_2175__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i29.GSR = "ENABLED";
    FD1S3IX count_2175__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i30.GSR = "ENABLED";
    FD1S3IX count_2175__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i31.GSR = "ENABLED";
    LUT4 i24683_2_lut (.A(n30948), .B(n34347), .Z(n2595)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24683_2_lut.init = 16'heeee;
    LUT4 i24681_4_lut (.A(n27), .B(n28180), .C(n25), .D(n26), .Z(n30948)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i24681_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n28180)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_374), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_431 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_431.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_432 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_432.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_374)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    CCU2D add_21615_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27952), 
          .S0(n6778));
    defparam add_21615_cout.INIT0 = 16'h0000;
    defparam add_21615_cout.INIT1 = 16'h0000;
    defparam add_21615_cout.INJECT1_0 = "NO";
    defparam add_21615_cout.INJECT1_1 = "NO";
    CCU2D add_21615_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27951), .COUT(n27952));
    defparam add_21615_24.INIT0 = 16'h5555;
    defparam add_21615_24.INIT1 = 16'h5555;
    defparam add_21615_24.INJECT1_0 = "NO";
    defparam add_21615_24.INJECT1_1 = "NO";
    CCU2D add_21615_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27950), .COUT(n27951));
    defparam add_21615_22.INIT0 = 16'h5555;
    defparam add_21615_22.INIT1 = 16'h5555;
    defparam add_21615_22.INJECT1_0 = "NO";
    defparam add_21615_22.INJECT1_1 = "NO";
    CCU2D add_21615_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27949), .COUT(n27950));
    defparam add_21615_20.INIT0 = 16'h5555;
    defparam add_21615_20.INIT1 = 16'h5555;
    defparam add_21615_20.INJECT1_0 = "NO";
    defparam add_21615_20.INJECT1_1 = "NO";
    CCU2D add_21615_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27948), .COUT(n27949));
    defparam add_21615_18.INIT0 = 16'h5555;
    defparam add_21615_18.INIT1 = 16'h5555;
    defparam add_21615_18.INJECT1_0 = "NO";
    defparam add_21615_18.INJECT1_1 = "NO";
    CCU2D add_21615_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27947), .COUT(n27948));
    defparam add_21615_16.INIT0 = 16'h5aaa;
    defparam add_21615_16.INIT1 = 16'h5555;
    defparam add_21615_16.INJECT1_0 = "NO";
    defparam add_21615_16.INJECT1_1 = "NO";
    CCU2D add_21615_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27946), .COUT(n27947));
    defparam add_21615_14.INIT0 = 16'h5aaa;
    defparam add_21615_14.INIT1 = 16'h5555;
    defparam add_21615_14.INJECT1_0 = "NO";
    defparam add_21615_14.INJECT1_1 = "NO";
    CCU2D add_21615_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27945), .COUT(n27946));
    defparam add_21615_12.INIT0 = 16'h5555;
    defparam add_21615_12.INIT1 = 16'h5aaa;
    defparam add_21615_12.INJECT1_0 = "NO";
    defparam add_21615_12.INJECT1_1 = "NO";
    CCU2D add_21615_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27944), .COUT(n27945));
    defparam add_21615_10.INIT0 = 16'h5aaa;
    defparam add_21615_10.INIT1 = 16'h5aaa;
    defparam add_21615_10.INJECT1_0 = "NO";
    defparam add_21615_10.INJECT1_1 = "NO";
    CCU2D add_21615_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27943), .COUT(n27944));
    defparam add_21615_8.INIT0 = 16'h5555;
    defparam add_21615_8.INIT1 = 16'h5aaa;
    defparam add_21615_8.INJECT1_0 = "NO";
    defparam add_21615_8.INJECT1_1 = "NO";
    CCU2D add_21615_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27942), .COUT(n27943));
    defparam add_21615_6.INIT0 = 16'h5555;
    defparam add_21615_6.INIT1 = 16'h5555;
    defparam add_21615_6.INJECT1_0 = "NO";
    defparam add_21615_6.INJECT1_1 = "NO";
    CCU2D add_21615_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27941), .COUT(n27942));
    defparam add_21615_4.INIT0 = 16'h5aaa;
    defparam add_21615_4.INIT1 = 16'h5aaa;
    defparam add_21615_4.INJECT1_0 = "NO";
    defparam add_21615_4.INJECT1_1 = "NO";
    CCU2D add_21615_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27941));
    defparam add_21615_2.INIT0 = 16'h7000;
    defparam add_21615_2.INIT1 = 16'h5555;
    defparam add_21615_2.INJECT1_0 = "NO";
    defparam add_21615_2.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27858), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_33.INIT1 = 16'h0000;
    defparam count_2175_add_4_33.INJECT1_0 = "NO";
    defparam count_2175_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27857), .COUT(n27858), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_31.INJECT1_0 = "NO";
    defparam count_2175_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27856), .COUT(n27857), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_29.INJECT1_0 = "NO";
    defparam count_2175_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27855), .COUT(n27856), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_27.INJECT1_0 = "NO";
    defparam count_2175_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27854), .COUT(n27855), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_25.INJECT1_0 = "NO";
    defparam count_2175_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27853), .COUT(n27854), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_23.INJECT1_0 = "NO";
    defparam count_2175_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27852), .COUT(n27853), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_21.INJECT1_0 = "NO";
    defparam count_2175_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27851), .COUT(n27852), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_19.INJECT1_0 = "NO";
    defparam count_2175_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27850), .COUT(n27851), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_17.INJECT1_0 = "NO";
    defparam count_2175_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27849), .COUT(n27850), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_15.INJECT1_0 = "NO";
    defparam count_2175_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27848), .COUT(n27849), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_13.INJECT1_0 = "NO";
    defparam count_2175_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27847), .COUT(n27848), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_11.INJECT1_0 = "NO";
    defparam count_2175_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27846), .COUT(n27847), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_9.INJECT1_0 = "NO";
    defparam count_2175_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27845), .COUT(n27846), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_7.INJECT1_0 = "NO";
    defparam count_2175_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27844), .COUT(n27845), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_5.INJECT1_0 = "NO";
    defparam count_2175_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27843), .COUT(n27844), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_3.INJECT1_0 = "NO";
    defparam count_2175_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27843), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_1.INIT0 = 16'hF000;
    defparam count_2175_add_4_1.INIT1 = 16'h0555;
    defparam count_2175_add_4_1.INJECT1_0 = "NO";
    defparam count_2175_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (n34344, n32422, \register_addr[5] , 
            n30431, read_value, debug_c_c, n11981, n32400, \register_addr[1] , 
            VCC_net, GND_net, Stepper_Z_nFault_c, n34349, \read_size[0] , 
            n30658, Stepper_Z_M0_c_0, n579, prev_select, n32449, n32534, 
            n32442, rw, n34347, n32396, n7852, n34350, databus, 
            n608, n610, \control_reg[7] , Stepper_Z_En_c, n34351, 
            Stepper_Z_Dir_c, Stepper_Z_M2_c_2, Stepper_Z_M1_c_1, \read_size[2] , 
            n29690, \steps_reg[5] , \steps_reg[3] , n34352, n14, \register_addr[0] , 
            n15, stepping, n30316, n32473, n32525, n32395, n20528, 
            limit_c_2, n28214, Stepper_Z_Step_c, n32463) /* synthesis syn_module_defined=1 */ ;
    input n34344;
    input n32422;
    input \register_addr[5] ;
    input n30431;
    output [31:0]read_value;
    input debug_c_c;
    input n11981;
    input n32400;
    input \register_addr[1] ;
    input VCC_net;
    input GND_net;
    input Stepper_Z_nFault_c;
    input n34349;
    output \read_size[0] ;
    input n30658;
    output Stepper_Z_M0_c_0;
    input n579;
    output prev_select;
    input n32449;
    input n32534;
    input n32442;
    input rw;
    input n34347;
    input n32396;
    input n7852;
    input n34350;
    input [31:0]databus;
    input n608;
    input n610;
    output \control_reg[7] ;
    output Stepper_Z_En_c;
    input n34351;
    output Stepper_Z_Dir_c;
    output Stepper_Z_M2_c_2;
    output Stepper_Z_M1_c_1;
    output \read_size[2] ;
    input n29690;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input n34352;
    input n14;
    input \register_addr[0] ;
    input n15;
    input stepping;
    input n30316;
    input n32473;
    input n32525;
    input n32395;
    output n20528;
    input limit_c_2;
    output n28214;
    output Stepper_Z_Step_c;
    input n32463;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n3276, n30843, n30886, n30887, n30888, fault_latched;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n3277;
    
    wire n12372, prev_step_clk, step_clk, limit_latched, n182, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n12358, n32381, n9610;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]n224;
    
    wire n30924;
    wire [31:0]n5782;
    
    wire n18868, n6;
    wire [7:0]n7333;
    wire [31:0]n5746;
    
    wire n30322, n30319, n30323, n30324, n30325, n30326, n30327, 
        n30328, n30329, n30330, n30331, n30320, n30332, n30333, 
        n30334, n30335, n30321, n30336, n30337, n30338, n30339, 
        n30340, n30317, n30318, int_step, n20522, n32394, n30922, 
        n30923, n18866, n18869, n5, n27754, n27753, n27752, n27751, 
        n27750, n30841, n30842, n27749, n27748, n27747, n27746, 
        n27745, n27744, n27743, n27742, n27741, n27740, n27739, 
        n49, n62, n58, n50, n41, n60, n54, n42, n52, n38, 
        n56, n46;
    
    LUT4 i2_3_lut_4_lut (.A(n34344), .B(n32422), .C(\register_addr[5] ), 
         .D(n30431), .Z(n3276)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_4_lut.init = 16'h4000;
    FD1P3IX read_value__i0 (.D(n30843), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    PFUMX i24530 (.BLUT(n30886), .ALUT(n30887), .C0(\register_addr[1] ), 
          .Z(n30888));
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3277[0]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n30658), .SP(n11981), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12372), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12358), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32449), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i24748_3_lut_rep_256_4_lut_4_lut (.A(n32534), .B(n32442), .C(n32422), 
         .D(rw), .Z(n32381)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24748_3_lut_rep_256_4_lut_4_lut.init = 16'h0010;
    LUT4 i24776_2_lut_4_lut_4_lut (.A(n32534), .B(n34347), .C(n32396), 
         .D(n32442), .Z(n12372)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24776_2_lut_4_lut_4_lut.init = 16'hccdc;
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n7852), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n7852), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n7852), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n7852), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n7852), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n7852), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n7852), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n12358), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12358), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n32381), .CD(n9610), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n32381), .PD(n34351), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n32381), .PD(n34351), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n12372), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n32381), .PD(n34351), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n12372), .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n32381), .PD(n34351), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n29690), .SP(n11981), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3277[31]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3277[30]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3277[29]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3277[28]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3277[27]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3277[26]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3277[25]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3277[24]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3277[23]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3277[22]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3277[21]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3277[20]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3277[19]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3277[18]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3277[17]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3277[16]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3277[15]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3277[14]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3277[13]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3277[12]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3277[11]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3277[10]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3277[9]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3277[8]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3277[7]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3277[6]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3277[5]), .CK(debug_c_c), .CD(n34351), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3277[4]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3277[3]), .CK(debug_c_c), .CD(n34352), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3277[2]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3277[1]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1338_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3276), 
         .Z(n3277[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i32_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i1 (.D(n30924), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1338_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3276), 
         .Z(n3277[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3276), 
         .Z(n3277[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3276), 
         .Z(n3277[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3276), 
         .Z(n3277[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3276), 
         .Z(n3277[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3276), 
         .Z(n3277[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3276), 
         .Z(n3277[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3276), 
         .Z(n3277[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3276), 
         .Z(n3277[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3276), 
         .Z(n3277[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3276), 
         .Z(n3277[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3276), 
         .Z(n3277[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3276), 
         .Z(n3277[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i19_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i2 (.D(n30888), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5782[3]), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5782[4]), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18868), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 mux_1338_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3276), 
         .Z(n3277[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i18_3_lut.init = 16'hcaca;
    PFUMX mux_1650_i5 (.BLUT(n7333[4]), .ALUT(n5746[4]), .C0(\register_addr[1] ), 
          .Z(n5782[4]));
    PFUMX mux_1650_i8 (.BLUT(n7333[7]), .ALUT(n5746[7]), .C0(\register_addr[1] ), 
          .Z(n5782[7]));
    FD1P3IX read_value__i7 (.D(n5782[7]), .SP(n11981), .CD(n32400), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30322), .SP(n11981), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n30319), .SP(n11981), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    LUT4 mux_1338_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3276), 
         .Z(n3277[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i17_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i10 (.D(n30323), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    LUT4 mux_1338_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3276), 
         .Z(n3277[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i16_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i11 (.D(n30324), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30325), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30326), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30327), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n30328), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n30329), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n30330), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n30331), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30320), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30332), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30333), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30334), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30335), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30321), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    LUT4 mux_1338_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3276), 
         .Z(n3277[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3276), 
         .Z(n3277[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3276), 
         .Z(n3277[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3276), 
         .Z(n3277[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3276), 
         .Z(n3277[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3276), .Z(n3277[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3276), .Z(n3277[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3276), .Z(n3277[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3276), .Z(n3277[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i7_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i25 (.D(n30336), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n30337), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30338), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30339), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30340), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30317), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n30318), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n32394), .SP(n20522), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1338_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3276), .Z(n3277[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3276), .Z(n3277[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3276), .Z(n3277[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3276), .Z(n3277[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3276), .Z(n3277[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i2_3_lut.init = 16'hcaca;
    LUT4 i24564_3_lut (.A(Stepper_Z_M1_c_1), .B(div_factor_reg[1]), .C(\register_addr[1] ), 
         .Z(n30922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24564_3_lut.init = 16'hcaca;
    LUT4 i24565_3_lut (.A(fault_latched), .B(steps_reg[1]), .C(\register_addr[1] ), 
         .Z(n30923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24565_3_lut.init = 16'hcaca;
    PFUMX i13127 (.BLUT(n18866), .ALUT(n14), .C0(\register_addr[0] ), 
          .Z(n18868));
    PFUMX i13130 (.BLUT(n18869), .ALUT(n15), .C0(\register_addr[0] ), 
          .Z(n5782[3]));
    PFUMX i6 (.BLUT(n7333[6]), .ALUT(n5), .C0(\register_addr[1] ), .Z(n6));
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27754), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    LUT4 i14008_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7333[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14008_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27753), .COUT(n27754), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27752), .COUT(n27753), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    LUT4 mux_1646_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5746[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1646_i5_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27751), .COUT(n27752), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    LUT4 mux_1338_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3276), .Z(n3277[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i1_3_lut.init = 16'hcaca;
    LUT4 i14006_2_lut (.A(\control_reg[7] ), .B(\register_addr[0] ), .Z(n7333[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14006_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27750), .COUT(n27751), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    PFUMX i24485 (.BLUT(n30841), .ALUT(n30842), .C0(\register_addr[1] ), 
          .Z(n30843));
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27749), .COUT(n27750), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27748), .COUT(n27749), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27747), .COUT(n27748), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27746), .COUT(n27747), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27745), .COUT(n27746), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27744), .COUT(n27745), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27743), .COUT(n27744), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27742), .COUT(n27743), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27741), .COUT(n27742), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27740), .COUT(n27741), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27739), .COUT(n27740), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27739), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_1646_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5746[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1646_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(div_factor_reg[8]), .B(n30316), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n30322)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_408 (.A(div_factor_reg[9]), .B(n30316), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n30319)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_408.init = 16'hc088;
    LUT4 i1_4_lut_adj_409 (.A(div_factor_reg[10]), .B(n30316), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n30323)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_409.init = 16'hc088;
    LUT4 i1_4_lut_adj_410 (.A(div_factor_reg[11]), .B(n30316), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n30324)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_410.init = 16'hc088;
    LUT4 i1_4_lut_adj_411 (.A(div_factor_reg[12]), .B(n30316), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n30325)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_411.init = 16'hc088;
    LUT4 i1_4_lut_adj_412 (.A(div_factor_reg[13]), .B(n30316), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n30326)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_412.init = 16'hc088;
    LUT4 i2_3_lut_rep_269 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n32394)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_269.init = 16'h0808;
    LUT4 i14784_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n34347), .Z(n20522)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14784_4_lut_4_lut.init = 16'h0038;
    LUT4 i24793_2_lut_3_lut_3_lut_4_lut (.A(n32473), .B(n32525), .C(n32395), 
         .D(n34347), .Z(n20528)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24793_2_lut_3_lut_3_lut_4_lut.init = 16'hff10;
    LUT4 i1_4_lut_adj_413 (.A(div_factor_reg[14]), .B(n30316), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n30327)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_413.init = 16'hc088;
    LUT4 i1_4_lut_adj_414 (.A(div_factor_reg[15]), .B(n30316), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n30328)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_414.init = 16'hc088;
    LUT4 i1_4_lut_adj_415 (.A(div_factor_reg[16]), .B(n30316), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n30329)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_415.init = 16'hc088;
    LUT4 i1_4_lut_adj_416 (.A(div_factor_reg[17]), .B(n30316), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n30330)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_416.init = 16'hc088;
    LUT4 i1_4_lut_adj_417 (.A(div_factor_reg[18]), .B(n30316), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n30331)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_417.init = 16'hc088;
    LUT4 i1_4_lut_adj_418 (.A(div_factor_reg[19]), .B(n30316), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n30320)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_418.init = 16'hc088;
    LUT4 i1_4_lut_adj_419 (.A(div_factor_reg[20]), .B(n30316), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n30332)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_419.init = 16'hc088;
    LUT4 i1_4_lut_adj_420 (.A(div_factor_reg[21]), .B(n30316), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n30333)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_420.init = 16'hc088;
    LUT4 i1_4_lut_adj_421 (.A(div_factor_reg[22]), .B(n30316), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n30334)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_421.init = 16'hc088;
    LUT4 i1_4_lut_adj_422 (.A(div_factor_reg[23]), .B(n30316), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n30335)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_422.init = 16'hc088;
    LUT4 i1_4_lut_adj_423 (.A(div_factor_reg[24]), .B(n30316), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n30321)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_423.init = 16'hc088;
    LUT4 i1_4_lut_adj_424 (.A(div_factor_reg[25]), .B(n30316), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n30336)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_424.init = 16'hc088;
    LUT4 i1_4_lut_adj_425 (.A(div_factor_reg[26]), .B(n30316), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n30337)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_425.init = 16'hc088;
    LUT4 i1_4_lut_adj_426 (.A(div_factor_reg[27]), .B(n30316), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n30338)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_426.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_427 (.A(div_factor_reg[28]), .B(n30316), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n30339)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_427.init = 16'hc088;
    LUT4 i1_2_lut (.A(n7852), .B(n34347), .Z(n12358)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_428 (.A(div_factor_reg[29]), .B(n30316), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n30340)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_428.init = 16'hc088;
    LUT4 i1_4_lut_adj_429 (.A(div_factor_reg[30]), .B(n30316), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n30317)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_429.init = 16'hc088;
    LUT4 i1_4_lut_adj_430 (.A(div_factor_reg[31]), .B(n30316), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n30318)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_430.init = 16'hc088;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12358), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i13125_3_lut (.A(Stepper_Z_Dir_c), .B(div_factor_reg[5]), .C(\register_addr[1] ), 
         .Z(n18866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13125_3_lut.init = 16'hcaca;
    LUT4 i13128_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(\register_addr[1] ), 
         .Z(n18869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13128_3_lut.init = 16'hcaca;
    LUT4 i14007_2_lut (.A(Stepper_Z_En_c), .B(\register_addr[0] ), .Z(n7333[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14007_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    LUT4 i24528_3_lut (.A(Stepper_Z_M2_c_2), .B(stepping), .C(\register_addr[0] ), 
         .Z(n30886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24528_3_lut.init = 16'hcaca;
    LUT4 i24529_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24529_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28214)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i24483_3_lut (.A(Stepper_Z_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24483_3_lut.init = 16'hcaca;
    LUT4 i17_4_lut (.A(steps_reg[24]), .B(steps_reg[20]), .C(steps_reg[9]), 
         .D(steps_reg[1]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i24484_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24484_3_lut.init = 16'hcaca;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[2]), .B(n52), .C(n38), .D(steps_reg[4]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[0]), .B(steps_reg[10]), .C(steps_reg[28]), 
         .D(\steps_reg[3] ), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[12]), .B(steps_reg[18]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[22]), .B(n56), .C(n46), .D(\steps_reg[5] ), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[30]), .B(steps_reg[14]), .C(steps_reg[7]), 
         .D(steps_reg[19]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i24669_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i24669_2_lut.init = 16'h9999;
    LUT4 i10_2_lut (.A(steps_reg[16]), .B(steps_reg[27]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[23]), .B(steps_reg[13]), .C(steps_reg[29]), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[17]), .B(steps_reg[15]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[21]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[8]), .B(steps_reg[11]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i6_2_lut.init = 16'heeee;
    PFUMX i24566 (.BLUT(n30922), .ALUT(n30923), .C0(\register_addr[0] ), 
          .Z(n30924));
    LUT4 i3849_3_lut (.A(prev_limit_latched), .B(n34347), .C(limit_latched), 
         .Z(n9610)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3849_3_lut.init = 16'hdcdc;
    ClockDivider step_clk_gen (.debug_c_c(debug_c_c), .div_factor_reg({div_factor_reg}), 
            .n34347(n34347), .step_clk(step_clk), .n32463(n32463), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (debug_c_c, div_factor_reg, n34347, step_clk, n32463, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input n34347;
    output step_clk;
    input n32463;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n32372, n14407, n7056, n7090, n7021;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27421;
    wire [31:0]n40;
    
    wire n27422, n27420, n27419, n27418, n27417, n27416, n27415, 
        n27414, n27413, n27412, n27411, n27410, n27409, n27690, 
        n27689, n27408, n27407, n27688, n27687, n27406, n27405, 
        n27686, n27685, n27404, n27684, n27683, n27403, n27402, 
        n27682, n27681, n27401, n27680, n27679, n27400, n27678, 
        n27399, n27677, n27398, n27397, n27676, n27396, n27675, 
        n27395, n27394, n27393, n27392, n27391, n27438, n27437, 
        n27436, n27435, n27434, n27433, n27432, n27431, n27430, 
        n27429, n27428, n27427, n27426, n27425, n27424, n27423, 
        n27810, n27809, n27808, n27807, n27806, n27805, n27804, 
        n27803, n27802, n27801, n27800, n27799, n27798, n27797, 
        n27796, n27795;
    
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    LUT4 i962_2_lut_rep_247 (.A(n7056), .B(n34347), .Z(n32372)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i962_2_lut_rep_247.init = 16'heeee;
    LUT4 i8641_2_lut_3_lut (.A(n7056), .B(n34347), .C(n7090), .Z(n14407)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8641_2_lut_3_lut.init = 16'he0e0;
    FD1S3IX clk_o_22 (.D(n7021), .CK(debug_c_c), .CD(n32463), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2178__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i0.GSR = "ENABLED";
    FD1S3IX count_2178__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i1.GSR = "ENABLED";
    FD1S3IX count_2178__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i2.GSR = "ENABLED";
    FD1S3IX count_2178__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i3.GSR = "ENABLED";
    FD1S3IX count_2178__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i4.GSR = "ENABLED";
    FD1S3IX count_2178__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i5.GSR = "ENABLED";
    FD1S3IX count_2178__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i6.GSR = "ENABLED";
    FD1S3IX count_2178__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i7.GSR = "ENABLED";
    FD1S3IX count_2178__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i8.GSR = "ENABLED";
    FD1S3IX count_2178__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i9.GSR = "ENABLED";
    FD1S3IX count_2178__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i10.GSR = "ENABLED";
    FD1S3IX count_2178__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i11.GSR = "ENABLED";
    FD1S3IX count_2178__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i12.GSR = "ENABLED";
    FD1S3IX count_2178__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i13.GSR = "ENABLED";
    FD1S3IX count_2178__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i14.GSR = "ENABLED";
    FD1S3IX count_2178__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i15.GSR = "ENABLED";
    FD1S3IX count_2178__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i16.GSR = "ENABLED";
    FD1S3IX count_2178__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i17.GSR = "ENABLED";
    FD1S3IX count_2178__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i18.GSR = "ENABLED";
    FD1S3IX count_2178__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i19.GSR = "ENABLED";
    FD1S3IX count_2178__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i20.GSR = "ENABLED";
    FD1S3IX count_2178__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i21.GSR = "ENABLED";
    FD1S3IX count_2178__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i22.GSR = "ENABLED";
    FD1S3IX count_2178__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i23.GSR = "ENABLED";
    FD1S3IX count_2178__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i24.GSR = "ENABLED";
    FD1S3IX count_2178__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i25.GSR = "ENABLED";
    FD1S3IX count_2178__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i26.GSR = "ENABLED";
    FD1S3IX count_2178__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i27.GSR = "ENABLED";
    FD1S3IX count_2178__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i28.GSR = "ENABLED";
    FD1S3IX count_2178__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i29.GSR = "ENABLED";
    FD1S3IX count_2178__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i30.GSR = "ENABLED";
    FD1S3IX count_2178__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32372), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    CCU2D sub_1726_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27421), .COUT(n27422));
    defparam sub_1726_add_2_31.INIT0 = 16'h5999;
    defparam sub_1726_add_2_31.INIT1 = 16'h5999;
    defparam sub_1726_add_2_31.INJECT1_0 = "NO";
    defparam sub_1726_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27420), .COUT(n27421));
    defparam sub_1726_add_2_29.INIT0 = 16'h5999;
    defparam sub_1726_add_2_29.INIT1 = 16'h5999;
    defparam sub_1726_add_2_29.INJECT1_0 = "NO";
    defparam sub_1726_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27419), .COUT(n27420));
    defparam sub_1726_add_2_27.INIT0 = 16'h5999;
    defparam sub_1726_add_2_27.INIT1 = 16'h5999;
    defparam sub_1726_add_2_27.INJECT1_0 = "NO";
    defparam sub_1726_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27418), .COUT(n27419));
    defparam sub_1726_add_2_25.INIT0 = 16'h5999;
    defparam sub_1726_add_2_25.INIT1 = 16'h5999;
    defparam sub_1726_add_2_25.INJECT1_0 = "NO";
    defparam sub_1726_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27417), .COUT(n27418));
    defparam sub_1726_add_2_23.INIT0 = 16'h5999;
    defparam sub_1726_add_2_23.INIT1 = 16'h5999;
    defparam sub_1726_add_2_23.INJECT1_0 = "NO";
    defparam sub_1726_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27416), .COUT(n27417));
    defparam sub_1726_add_2_21.INIT0 = 16'h5999;
    defparam sub_1726_add_2_21.INIT1 = 16'h5999;
    defparam sub_1726_add_2_21.INJECT1_0 = "NO";
    defparam sub_1726_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27415), .COUT(n27416));
    defparam sub_1726_add_2_19.INIT0 = 16'h5999;
    defparam sub_1726_add_2_19.INIT1 = 16'h5999;
    defparam sub_1726_add_2_19.INJECT1_0 = "NO";
    defparam sub_1726_add_2_19.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    CCU2D sub_1726_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27414), .COUT(n27415));
    defparam sub_1726_add_2_17.INIT0 = 16'h5999;
    defparam sub_1726_add_2_17.INIT1 = 16'h5999;
    defparam sub_1726_add_2_17.INJECT1_0 = "NO";
    defparam sub_1726_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27413), .COUT(n27414));
    defparam sub_1726_add_2_15.INIT0 = 16'h5999;
    defparam sub_1726_add_2_15.INIT1 = 16'h5999;
    defparam sub_1726_add_2_15.INJECT1_0 = "NO";
    defparam sub_1726_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27412), .COUT(n27413));
    defparam sub_1726_add_2_13.INIT0 = 16'h5999;
    defparam sub_1726_add_2_13.INIT1 = 16'h5999;
    defparam sub_1726_add_2_13.INJECT1_0 = "NO";
    defparam sub_1726_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27411), .COUT(n27412));
    defparam sub_1726_add_2_11.INIT0 = 16'h5999;
    defparam sub_1726_add_2_11.INIT1 = 16'h5999;
    defparam sub_1726_add_2_11.INJECT1_0 = "NO";
    defparam sub_1726_add_2_11.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    CCU2D sub_1726_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27410), .COUT(n27411));
    defparam sub_1726_add_2_9.INIT0 = 16'h5999;
    defparam sub_1726_add_2_9.INIT1 = 16'h5999;
    defparam sub_1726_add_2_9.INJECT1_0 = "NO";
    defparam sub_1726_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27409), .COUT(n27410));
    defparam sub_1726_add_2_7.INIT0 = 16'h5999;
    defparam sub_1726_add_2_7.INIT1 = 16'h5999;
    defparam sub_1726_add_2_7.INJECT1_0 = "NO";
    defparam sub_1726_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27690), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27689), .COUT(n27690), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27408), .COUT(n27409));
    defparam sub_1726_add_2_5.INIT0 = 16'h5999;
    defparam sub_1726_add_2_5.INIT1 = 16'h5999;
    defparam sub_1726_add_2_5.INJECT1_0 = "NO";
    defparam sub_1726_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27407), .COUT(n27408));
    defparam sub_1726_add_2_3.INIT0 = 16'h5999;
    defparam sub_1726_add_2_3.INIT1 = 16'h5999;
    defparam sub_1726_add_2_3.INJECT1_0 = "NO";
    defparam sub_1726_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32372), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27688), .COUT(n27689), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27407));
    defparam sub_1726_add_2_1.INIT0 = 16'h0000;
    defparam sub_1726_add_2_1.INIT1 = 16'h5999;
    defparam sub_1726_add_2_1.INJECT1_0 = "NO";
    defparam sub_1726_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27687), .COUT(n27688), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32372), .PD(n14407), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_1727_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27406), .S1(n7090));
    defparam sub_1727_add_2_33.INIT0 = 16'hf555;
    defparam sub_1727_add_2_33.INIT1 = 16'h0000;
    defparam sub_1727_add_2_33.INJECT1_0 = "NO";
    defparam sub_1727_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27405), .COUT(n27406));
    defparam sub_1727_add_2_31.INIT0 = 16'hf555;
    defparam sub_1727_add_2_31.INIT1 = 16'hf555;
    defparam sub_1727_add_2_31.INJECT1_0 = "NO";
    defparam sub_1727_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27686), .COUT(n27687), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27685), .COUT(n27686), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27404), .COUT(n27405));
    defparam sub_1727_add_2_29.INIT0 = 16'hf555;
    defparam sub_1727_add_2_29.INIT1 = 16'hf555;
    defparam sub_1727_add_2_29.INJECT1_0 = "NO";
    defparam sub_1727_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27684), .COUT(n27685), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27683), .COUT(n27684), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27403), .COUT(n27404));
    defparam sub_1727_add_2_27.INIT0 = 16'hf555;
    defparam sub_1727_add_2_27.INIT1 = 16'hf555;
    defparam sub_1727_add_2_27.INJECT1_0 = "NO";
    defparam sub_1727_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27402), .COUT(n27403));
    defparam sub_1727_add_2_25.INIT0 = 16'hf555;
    defparam sub_1727_add_2_25.INIT1 = 16'hf555;
    defparam sub_1727_add_2_25.INJECT1_0 = "NO";
    defparam sub_1727_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27682), .COUT(n27683), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27681), .COUT(n27682), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27401), .COUT(n27402));
    defparam sub_1727_add_2_23.INIT0 = 16'hf555;
    defparam sub_1727_add_2_23.INIT1 = 16'hf555;
    defparam sub_1727_add_2_23.INJECT1_0 = "NO";
    defparam sub_1727_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27680), .COUT(n27681), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27679), .COUT(n27680), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27400), .COUT(n27401));
    defparam sub_1727_add_2_21.INIT0 = 16'hf555;
    defparam sub_1727_add_2_21.INIT1 = 16'hf555;
    defparam sub_1727_add_2_21.INJECT1_0 = "NO";
    defparam sub_1727_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27678), .COUT(n27679), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27399), .COUT(n27400));
    defparam sub_1727_add_2_19.INIT0 = 16'hf555;
    defparam sub_1727_add_2_19.INIT1 = 16'hf555;
    defparam sub_1727_add_2_19.INJECT1_0 = "NO";
    defparam sub_1727_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27677), .COUT(n27678), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27398), .COUT(n27399));
    defparam sub_1727_add_2_17.INIT0 = 16'hf555;
    defparam sub_1727_add_2_17.INIT1 = 16'hf555;
    defparam sub_1727_add_2_17.INJECT1_0 = "NO";
    defparam sub_1727_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27397), .COUT(n27398));
    defparam sub_1727_add_2_15.INIT0 = 16'hf555;
    defparam sub_1727_add_2_15.INIT1 = 16'hf555;
    defparam sub_1727_add_2_15.INJECT1_0 = "NO";
    defparam sub_1727_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27676), .COUT(n27677), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27396), .COUT(n27397));
    defparam sub_1727_add_2_13.INIT0 = 16'hf555;
    defparam sub_1727_add_2_13.INIT1 = 16'hf555;
    defparam sub_1727_add_2_13.INJECT1_0 = "NO";
    defparam sub_1727_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27675), .COUT(n27676), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27395), .COUT(n27396));
    defparam sub_1727_add_2_11.INIT0 = 16'hf555;
    defparam sub_1727_add_2_11.INIT1 = 16'hf555;
    defparam sub_1727_add_2_11.INJECT1_0 = "NO";
    defparam sub_1727_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27394), .COUT(n27395));
    defparam sub_1727_add_2_9.INIT0 = 16'hf555;
    defparam sub_1727_add_2_9.INIT1 = 16'hf555;
    defparam sub_1727_add_2_9.INJECT1_0 = "NO";
    defparam sub_1727_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27675), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27393), .COUT(n27394));
    defparam sub_1727_add_2_7.INIT0 = 16'hf555;
    defparam sub_1727_add_2_7.INIT1 = 16'hf555;
    defparam sub_1727_add_2_7.INJECT1_0 = "NO";
    defparam sub_1727_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27392), .COUT(n27393));
    defparam sub_1727_add_2_5.INIT0 = 16'hf555;
    defparam sub_1727_add_2_5.INIT1 = 16'hf555;
    defparam sub_1727_add_2_5.INJECT1_0 = "NO";
    defparam sub_1727_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27391), .COUT(n27392));
    defparam sub_1727_add_2_3.INIT0 = 16'hf555;
    defparam sub_1727_add_2_3.INIT1 = 16'hf555;
    defparam sub_1727_add_2_3.INJECT1_0 = "NO";
    defparam sub_1727_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27391));
    defparam sub_1727_add_2_1.INIT0 = 16'h0000;
    defparam sub_1727_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1727_add_2_1.INJECT1_0 = "NO";
    defparam sub_1727_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27438), .S1(n7021));
    defparam sub_1724_add_2_33.INIT0 = 16'h5555;
    defparam sub_1724_add_2_33.INIT1 = 16'h0000;
    defparam sub_1724_add_2_33.INJECT1_0 = "NO";
    defparam sub_1724_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27437), .COUT(n27438));
    defparam sub_1724_add_2_31.INIT0 = 16'h5999;
    defparam sub_1724_add_2_31.INIT1 = 16'h5999;
    defparam sub_1724_add_2_31.INJECT1_0 = "NO";
    defparam sub_1724_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27436), .COUT(n27437));
    defparam sub_1724_add_2_29.INIT0 = 16'h5999;
    defparam sub_1724_add_2_29.INIT1 = 16'h5999;
    defparam sub_1724_add_2_29.INJECT1_0 = "NO";
    defparam sub_1724_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27435), .COUT(n27436));
    defparam sub_1724_add_2_27.INIT0 = 16'h5999;
    defparam sub_1724_add_2_27.INIT1 = 16'h5999;
    defparam sub_1724_add_2_27.INJECT1_0 = "NO";
    defparam sub_1724_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27434), .COUT(n27435));
    defparam sub_1724_add_2_25.INIT0 = 16'h5999;
    defparam sub_1724_add_2_25.INIT1 = 16'h5999;
    defparam sub_1724_add_2_25.INJECT1_0 = "NO";
    defparam sub_1724_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27433), .COUT(n27434));
    defparam sub_1724_add_2_23.INIT0 = 16'h5999;
    defparam sub_1724_add_2_23.INIT1 = 16'h5999;
    defparam sub_1724_add_2_23.INJECT1_0 = "NO";
    defparam sub_1724_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27432), .COUT(n27433));
    defparam sub_1724_add_2_21.INIT0 = 16'h5999;
    defparam sub_1724_add_2_21.INIT1 = 16'h5999;
    defparam sub_1724_add_2_21.INJECT1_0 = "NO";
    defparam sub_1724_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27431), .COUT(n27432));
    defparam sub_1724_add_2_19.INIT0 = 16'h5999;
    defparam sub_1724_add_2_19.INIT1 = 16'h5999;
    defparam sub_1724_add_2_19.INJECT1_0 = "NO";
    defparam sub_1724_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27430), .COUT(n27431));
    defparam sub_1724_add_2_17.INIT0 = 16'h5999;
    defparam sub_1724_add_2_17.INIT1 = 16'h5999;
    defparam sub_1724_add_2_17.INJECT1_0 = "NO";
    defparam sub_1724_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27429), .COUT(n27430));
    defparam sub_1724_add_2_15.INIT0 = 16'h5999;
    defparam sub_1724_add_2_15.INIT1 = 16'h5999;
    defparam sub_1724_add_2_15.INJECT1_0 = "NO";
    defparam sub_1724_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27428), .COUT(n27429));
    defparam sub_1724_add_2_13.INIT0 = 16'h5999;
    defparam sub_1724_add_2_13.INIT1 = 16'h5999;
    defparam sub_1724_add_2_13.INJECT1_0 = "NO";
    defparam sub_1724_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27427), .COUT(n27428));
    defparam sub_1724_add_2_11.INIT0 = 16'h5999;
    defparam sub_1724_add_2_11.INIT1 = 16'h5999;
    defparam sub_1724_add_2_11.INJECT1_0 = "NO";
    defparam sub_1724_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27426), .COUT(n27427));
    defparam sub_1724_add_2_9.INIT0 = 16'h5999;
    defparam sub_1724_add_2_9.INIT1 = 16'h5999;
    defparam sub_1724_add_2_9.INJECT1_0 = "NO";
    defparam sub_1724_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27425), .COUT(n27426));
    defparam sub_1724_add_2_7.INIT0 = 16'h5999;
    defparam sub_1724_add_2_7.INIT1 = 16'h5999;
    defparam sub_1724_add_2_7.INJECT1_0 = "NO";
    defparam sub_1724_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27424), .COUT(n27425));
    defparam sub_1724_add_2_5.INIT0 = 16'h5999;
    defparam sub_1724_add_2_5.INIT1 = 16'h5999;
    defparam sub_1724_add_2_5.INJECT1_0 = "NO";
    defparam sub_1724_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27423), .COUT(n27424));
    defparam sub_1724_add_2_3.INIT0 = 16'h5999;
    defparam sub_1724_add_2_3.INIT1 = 16'h5999;
    defparam sub_1724_add_2_3.INJECT1_0 = "NO";
    defparam sub_1724_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27423));
    defparam sub_1724_add_2_1.INIT0 = 16'h0000;
    defparam sub_1724_add_2_1.INIT1 = 16'h5999;
    defparam sub_1724_add_2_1.INJECT1_0 = "NO";
    defparam sub_1724_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27422), .S1(n7056));
    defparam sub_1726_add_2_33.INIT0 = 16'h5999;
    defparam sub_1726_add_2_33.INIT1 = 16'h0000;
    defparam sub_1726_add_2_33.INJECT1_0 = "NO";
    defparam sub_1726_add_2_33.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27810), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_33.INIT1 = 16'h0000;
    defparam count_2178_add_4_33.INJECT1_0 = "NO";
    defparam count_2178_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27809), .COUT(n27810), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_31.INJECT1_0 = "NO";
    defparam count_2178_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27808), .COUT(n27809), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_29.INJECT1_0 = "NO";
    defparam count_2178_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27807), .COUT(n27808), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_27.INJECT1_0 = "NO";
    defparam count_2178_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27806), .COUT(n27807), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_25.INJECT1_0 = "NO";
    defparam count_2178_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27805), .COUT(n27806), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_23.INJECT1_0 = "NO";
    defparam count_2178_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27804), .COUT(n27805), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_21.INJECT1_0 = "NO";
    defparam count_2178_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27803), .COUT(n27804), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_19.INJECT1_0 = "NO";
    defparam count_2178_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27802), .COUT(n27803), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_17.INJECT1_0 = "NO";
    defparam count_2178_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27801), .COUT(n27802), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_15.INJECT1_0 = "NO";
    defparam count_2178_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27800), .COUT(n27801), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_13.INJECT1_0 = "NO";
    defparam count_2178_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27799), .COUT(n27800), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_11.INJECT1_0 = "NO";
    defparam count_2178_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27798), .COUT(n27799), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_9.INJECT1_0 = "NO";
    defparam count_2178_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27797), .COUT(n27798), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_7.INJECT1_0 = "NO";
    defparam count_2178_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27796), .COUT(n27797), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_5.INJECT1_0 = "NO";
    defparam count_2178_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27795), .COUT(n27796), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_3.INJECT1_0 = "NO";
    defparam count_2178_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27795), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_1.INIT0 = 16'hF000;
    defparam count_2178_add_4_1.INIT1 = 16'h0555;
    defparam count_2178_add_4_1.INJECT1_0 = "NO";
    defparam count_2178_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (register_addr, read_value, 
            debug_c_c, n12620, GND_net, n34350, n3181, VCC_net, 
            Stepper_A_nFault_c, \read_size[0] , n30435, n32527, n32525, 
            n30311, Stepper_A_M0_c_0, n20528, n579, n12224, prev_select, 
            n32441, n32379, n34348, \databus[31] , \databus[28] , 
            n34349, \databus[13] , \databus[11] , \databus[10] , \databus[9] , 
            \databus[7] , \databus[6] , \databus[5] , n610, \control_reg[7] , 
            Stepper_A_En_c, Stepper_A_Dir_c, \databus[4] , \databus[3] , 
            Stepper_A_M2_c_2, Stepper_A_M1_c_1, \databus[1] , \read_size[2] , 
            n30363, n32396, n7852, n34351, n34352, \steps_reg[5] , 
            \steps_reg[3] , n32442, n32508, n32509, n32471, n14, 
            n15, n224, n32482, \register[2][0] , n15_adj_187, \register[2][3] , 
            n4, n32488, n32473, stepping, n34347, \databus[8] , 
            \databus[12] , \databus[14] , \databus[15] , \databus[16] , 
            \databus[17] , \databus[18] , \databus[19] , \databus[20] , 
            \databus[21] , \databus[22] , \databus[23] , \databus[24] , 
            \databus[25] , \databus[26] , \databus[27] , \databus[29] , 
            \databus[30] , limit_c_3, n32416, n30454, rw, n28299, 
            Stepper_A_Step_c, n32463) /* synthesis syn_module_defined=1 */ ;
    input [7:0]register_addr;
    output [31:0]read_value;
    input debug_c_c;
    input n12620;
    input GND_net;
    input n34350;
    input [31:0]n3181;
    input VCC_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n30435;
    output n32527;
    input n32525;
    output n30311;
    output Stepper_A_M0_c_0;
    input n20528;
    input n579;
    input n12224;
    output prev_select;
    input n32441;
    input n32379;
    input n34348;
    input \databus[31] ;
    input \databus[28] ;
    input n34349;
    input \databus[13] ;
    input \databus[11] ;
    input \databus[10] ;
    input \databus[9] ;
    input \databus[7] ;
    input \databus[6] ;
    input \databus[5] ;
    input n610;
    output \control_reg[7] ;
    output Stepper_A_En_c;
    output Stepper_A_Dir_c;
    input \databus[4] ;
    input \databus[3] ;
    output Stepper_A_M2_c_2;
    output Stepper_A_M1_c_1;
    input \databus[1] ;
    output \read_size[2] ;
    input n30363;
    input n32396;
    output n7852;
    input n34351;
    input n34352;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    output n32442;
    input n32508;
    input n32509;
    output n32471;
    input n14;
    input n15;
    output [31:0]n224;
    output n32482;
    input \register[2][0] ;
    output n15_adj_187;
    input \register[2][3] ;
    output n4;
    output n32488;
    output n32473;
    input stepping;
    input n34347;
    input \databus[8] ;
    input \databus[12] ;
    input \databus[14] ;
    input \databus[15] ;
    input \databus[16] ;
    input \databus[17] ;
    input \databus[18] ;
    input \databus[19] ;
    input \databus[20] ;
    input \databus[21] ;
    input \databus[22] ;
    input \databus[23] ;
    input \databus[24] ;
    input \databus[25] ;
    input \databus[26] ;
    input \databus[27] ;
    input \databus[29] ;
    input \databus[30] ;
    input limit_c_3;
    input n32416;
    input n30454;
    input rw;
    output n28299;
    output Stepper_A_Step_c;
    input n32463;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30892, n30893, n30894, n30846;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n56, n46, n60, fault_latched, prev_step_clk, step_clk, 
        limit_latched, n182, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n32380, n9608;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [7:0]n7342;
    wire [31:0]n6060;
    wire [31:0]n6096;
    
    wire n5, n6, int_step, n20536, n32392, n30855, n18830, n30401, 
        n30398, n30399, n30400, n30396;
    wire [31:0]n100;
    
    wire n30395, n30397, n30394, n30402, n30403, n30404, n30405, 
        n30406, n30407, n30408, n30409, n30410, n30411, n30412, 
        n30853, n30854, n30393, n18828, n18831, n30844, n30845, 
        n27738, n27737, n27736, n27735, n27734, n27733, n27732, 
        n27731, n27730, n27729, n54, n27728, n42, n27727, n27726, 
        n27725, n27724, n27723, n52, n38, n49, n62_adj_373, n58, 
        n50, n41;
    
    PFUMX i24536 (.BLUT(n30892), .ALUT(n30893), .C0(register_addr[1]), 
          .Z(n30894));
    FD1P3IX read_value__i0 (.D(n30846), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i28_4_lut (.A(steps_reg[20]), .B(n56), .C(n46), .D(steps_reg[15]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    FD1S3IX steps_reg__i0 (.D(n3181[0]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n30435), .SP(n12620), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(register_addr[5]), .B(register_addr[4]), .C(n32527), 
         .D(n32525), .Z(n30311)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0002;
    LUT4 equal_1407_i11_2_lut_rep_402 (.A(register_addr[2]), .B(register_addr[3]), 
         .Z(n32527)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_1407_i11_2_lut_rep_402.init = 16'heeee;
    FD1P3AX control_reg_i1 (.D(n579), .SP(n20528), .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12224), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32441), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(\databus[31] ), .SP(n32379), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(\databus[28] ), .SP(n32379), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(\databus[13] ), .SP(n32379), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(\databus[11] ), .SP(n32379), .PD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(\databus[10] ), .SP(n32379), .PD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(\databus[9] ), .SP(n32379), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(\databus[7] ), .SP(n32379), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(\databus[6] ), .SP(n32379), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(\databus[5] ), .SP(n32379), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12224), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(\databus[7] ), .SP(n32380), .CD(n9608), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(\databus[6] ), .SP(n32380), .PD(n34350), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(\databus[5] ), .SP(n32380), .PD(n34350), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(\databus[4] ), .SP(n32380), .CD(n34350), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(\databus[3] ), .SP(n32380), .PD(n34350), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n20528), .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(\databus[1] ), .SP(n32380), .PD(n34350), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n30363), .SP(n12620), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i3_4_lut_4_lut (.A(register_addr[1]), .B(register_addr[0]), .C(n32396), 
         .D(n30311), .Z(n7852)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i3_4_lut_4_lut.init = 16'h2000;
    FD1S3IX steps_reg__i31 (.D(n3181[31]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3181[30]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3181[29]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3181[28]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3181[27]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3181[26]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3181[25]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3181[24]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3181[23]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3181[22]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3181[21]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3181[20]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3181[19]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3181[18]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3181[17]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3181[16]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3181[15]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3181[14]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3181[13]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3181[12]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3181[11]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3181[10]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3181[9]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3181[8]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3181[7]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3181[6]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3181[5]), .CK(debug_c_c), .CD(n34352), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3181[4]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3181[3]), .CK(debug_c_c), .CD(n34352), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3181[2]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3181[1]), .CK(debug_c_c), .CD(n34352), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_317_3_lut_4_lut (.A(register_addr[1]), .B(n32527), 
         .C(n32525), .D(register_addr[0]), .Z(n32442)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(85[9:13])
    defparam i1_2_lut_rep_317_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_346_3_lut_4_lut (.A(register_addr[1]), .B(n32527), 
         .C(n32508), .D(n32509), .Z(n32471)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(85[9:13])
    defparam i1_2_lut_rep_346_3_lut_4_lut.init = 16'hfffe;
    PFUMX mux_1676_i5 (.BLUT(n7342[4]), .ALUT(n6060[4]), .C0(register_addr[1]), 
          .Z(n6096[4]));
    PFUMX mux_1676_i8 (.BLUT(n7342[7]), .ALUT(n6060[7]), .C0(register_addr[1]), 
          .Z(n6096[7]));
    PFUMX i6 (.BLUT(n7342[6]), .ALUT(n5), .C0(register_addr[1]), .Z(n6));
    FD1P3AX int_step_182 (.D(n32392), .SP(n20536), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30855), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30894), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6096[3]), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6096[4]), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18830), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6096[7]), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30401), .SP(n12620), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n30398), .SP(n12620), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n30399), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n30400), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30396), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n12620), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n12620), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n12620), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n12620), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30395), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30397), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30394), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30402), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30403), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30404), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30405), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30406), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n30407), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n30408), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30409), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30410), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30411), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30412), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    PFUMX i24497 (.BLUT(n30853), .ALUT(n30854), .C0(register_addr[1]), 
          .Z(n30855));
    FD1P3AX read_value__i31 (.D(n30393), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    PFUMX i13088 (.BLUT(n18828), .ALUT(n14), .C0(register_addr[0]), .Z(n18830));
    PFUMX i13091 (.BLUT(n18831), .ALUT(n15), .C0(register_addr[0]), .Z(n6096[3]));
    PFUMX i24488 (.BLUT(n30844), .ALUT(n30845), .C0(register_addr[1]), 
          .Z(n30846));
    LUT4 i13998_2_lut (.A(control_reg[4]), .B(register_addr[0]), .Z(n7342[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13998_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27738), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27737), .COUT(n27738), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    LUT4 i14577_2_lut_rep_357_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[6]), .D(register_addr[7]), .Z(n32482)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i14577_2_lut_rep_357_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1672_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(register_addr[0]), 
         .Z(n6060[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1672_i5_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut (.A(register_addr[2]), .B(register_addr[3]), .C(\register[2][0] ), 
         .Z(n15_adj_187)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_388 (.A(register_addr[2]), .B(register_addr[3]), 
         .C(\register[2][3] ), .Z(n4)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut_adj_388.init = 16'h1010;
    LUT4 i1_2_lut_rep_363_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .Z(n32488)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_363_3_lut.init = 16'hfefe;
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27736), .COUT(n27737), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27735), .COUT(n27736), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27734), .COUT(n27735), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_348_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n32473)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_348_3_lut_4_lut.init = 16'hfffe;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27733), .COUT(n27734), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27732), .COUT(n27733), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_267 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n32392)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_267.init = 16'h0808;
    LUT4 i14798_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n34347), .Z(n20536)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14798_4_lut_4_lut.init = 16'h0038;
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27731), .COUT(n27732), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27730), .COUT(n27731), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27729), .COUT(n27730), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[12]), .C(steps_reg[6]), 
         .D(steps_reg[18]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27728), .COUT(n27729), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27727), .COUT(n27728), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27726), .COUT(n27727), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27725), .COUT(n27726), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27724), .COUT(n27725), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27723), .COUT(n27724), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    LUT4 i24_4_lut (.A(steps_reg[13]), .B(steps_reg[17]), .C(\steps_reg[5] ), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i13996_2_lut (.A(\control_reg[7] ), .B(register_addr[0]), .Z(n7342[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13996_2_lut.init = 16'h2222;
    LUT4 mux_1672_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(register_addr[0]), 
         .Z(n6060[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1672_i8_3_lut.init = 16'hcaca;
    LUT4 i14_2_lut (.A(steps_reg[23]), .B(steps_reg[29]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27723), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i13997_2_lut (.A(Stepper_A_En_c), .B(register_addr[0]), .Z(n7342[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13997_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(register_addr[0]), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(div_factor_reg[8]), .B(register_addr[1]), .C(steps_reg[8]), 
         .D(register_addr[0]), .Z(n30401)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_389 (.A(div_factor_reg[9]), .B(register_addr[1]), 
         .C(steps_reg[9]), .D(register_addr[0]), .Z(n30398)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_389.init = 16'hc088;
    LUT4 i1_4_lut_adj_390 (.A(div_factor_reg[10]), .B(register_addr[1]), 
         .C(steps_reg[10]), .D(register_addr[0]), .Z(n30399)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_390.init = 16'hc088;
    LUT4 i1_4_lut_adj_391 (.A(div_factor_reg[11]), .B(register_addr[1]), 
         .C(steps_reg[11]), .D(register_addr[0]), .Z(n30400)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_391.init = 16'hc088;
    LUT4 i1_4_lut_adj_392 (.A(div_factor_reg[12]), .B(register_addr[1]), 
         .C(steps_reg[12]), .D(register_addr[0]), .Z(n30396)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_392.init = 16'hc088;
    LUT4 i13992_4_lut (.A(div_factor_reg[18]), .B(register_addr[1]), .C(steps_reg[18]), 
         .D(register_addr[0]), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13992_4_lut.init = 16'hc088;
    LUT4 i13993_4_lut (.A(div_factor_reg[17]), .B(register_addr[1]), .C(steps_reg[17]), 
         .D(register_addr[0]), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13993_4_lut.init = 16'hc088;
    LUT4 i13994_4_lut (.A(div_factor_reg[16]), .B(register_addr[1]), .C(steps_reg[16]), 
         .D(register_addr[0]), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13994_4_lut.init = 16'hc088;
    LUT4 i13995_4_lut (.A(div_factor_reg[15]), .B(register_addr[1]), .C(steps_reg[15]), 
         .D(register_addr[0]), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13995_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_393 (.A(div_factor_reg[13]), .B(register_addr[1]), 
         .C(steps_reg[13]), .D(register_addr[0]), .Z(n30395)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_393.init = 16'hc088;
    LUT4 i1_4_lut_adj_394 (.A(div_factor_reg[14]), .B(register_addr[1]), 
         .C(steps_reg[14]), .D(register_addr[0]), .Z(n30397)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_394.init = 16'hc088;
    LUT4 i1_4_lut_adj_395 (.A(div_factor_reg[19]), .B(register_addr[1]), 
         .C(steps_reg[19]), .D(register_addr[0]), .Z(n30394)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_395.init = 16'hc088;
    LUT4 i1_4_lut_adj_396 (.A(div_factor_reg[20]), .B(register_addr[1]), 
         .C(steps_reg[20]), .D(register_addr[0]), .Z(n30402)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_396.init = 16'hc088;
    LUT4 i1_4_lut_adj_397 (.A(div_factor_reg[21]), .B(register_addr[1]), 
         .C(steps_reg[21]), .D(register_addr[0]), .Z(n30403)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_397.init = 16'hc088;
    LUT4 i1_4_lut_adj_398 (.A(div_factor_reg[22]), .B(register_addr[1]), 
         .C(steps_reg[22]), .D(register_addr[0]), .Z(n30404)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_398.init = 16'hc088;
    LUT4 i1_4_lut_adj_399 (.A(div_factor_reg[23]), .B(register_addr[1]), 
         .C(steps_reg[23]), .D(register_addr[0]), .Z(n30405)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_399.init = 16'hc088;
    LUT4 i1_4_lut_adj_400 (.A(div_factor_reg[24]), .B(register_addr[1]), 
         .C(steps_reg[24]), .D(register_addr[0]), .Z(n30406)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_400.init = 16'hc088;
    LUT4 i24534_3_lut (.A(Stepper_A_M2_c_2), .B(stepping), .C(register_addr[0]), 
         .Z(n30892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24534_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_401 (.A(div_factor_reg[25]), .B(register_addr[1]), 
         .C(steps_reg[25]), .D(register_addr[0]), .Z(n30407)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_401.init = 16'hc088;
    FD1P3IX div_factor_reg_i1 (.D(\databus[1] ), .SP(n12224), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(\databus[3] ), .SP(n12224), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(\databus[4] ), .SP(n12224), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(\databus[8] ), .SP(n12224), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(\databus[12] ), .SP(n12224), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(\databus[14] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(\databus[15] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(\databus[16] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(\databus[17] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(\databus[18] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(\databus[19] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(\databus[20] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(\databus[21] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(\databus[22] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(\databus[23] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(\databus[24] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(\databus[25] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(\databus[26] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(\databus[27] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(\databus[29] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(\databus[30] ), .SP(n12224), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_402 (.A(div_factor_reg[26]), .B(register_addr[1]), 
         .C(steps_reg[26]), .D(register_addr[0]), .Z(n30408)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_402.init = 16'hc088;
    LUT4 i1_4_lut_adj_403 (.A(div_factor_reg[27]), .B(register_addr[1]), 
         .C(steps_reg[27]), .D(register_addr[0]), .Z(n30409)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_403.init = 16'hc088;
    LUT4 i20_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_404 (.A(div_factor_reg[28]), .B(register_addr[1]), 
         .C(steps_reg[28]), .D(register_addr[0]), .Z(n30410)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_404.init = 16'hc088;
    LUT4 i24535_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(register_addr[0]), 
         .Z(n30893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24535_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_405 (.A(div_factor_reg[29]), .B(register_addr[1]), 
         .C(steps_reg[29]), .D(register_addr[0]), .Z(n30411)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_405.init = 16'hc088;
    LUT4 i1_4_lut_adj_406 (.A(div_factor_reg[30]), .B(register_addr[1]), 
         .C(steps_reg[30]), .D(register_addr[0]), .Z(n30412)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_406.init = 16'hc088;
    LUT4 i24495_3_lut (.A(Stepper_A_M1_c_1), .B(fault_latched), .C(register_addr[0]), 
         .Z(n30853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24495_3_lut.init = 16'hcaca;
    LUT4 i24496_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(register_addr[0]), 
         .Z(n30854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24496_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_407 (.A(div_factor_reg[31]), .B(register_addr[1]), 
         .C(steps_reg[31]), .D(register_addr[0]), .Z(n30393)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_407.init = 16'hc088;
    LUT4 i24729_2_lut_rep_255_4_lut_4_lut (.A(n32442), .B(n32416), .C(n30454), 
         .D(rw), .Z(n32380)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24729_2_lut_rep_255_4_lut_4_lut.init = 16'h0040;
    LUT4 i6_2_lut (.A(steps_reg[10]), .B(\steps_reg[3] ), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i13086_3_lut (.A(Stepper_A_Dir_c), .B(div_factor_reg[5]), .C(register_addr[1]), 
         .Z(n18828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13086_3_lut.init = 16'hcaca;
    LUT4 i13089_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(register_addr[1]), 
         .Z(n18831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13089_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_373), .C(n58), .D(n50), .Z(n28299)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg[9]), .C(steps_reg[28]), 
         .D(steps_reg[2]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i24486_3_lut (.A(Stepper_A_M0_c_0), .B(limit_latched), .C(register_addr[0]), 
         .Z(n30844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24486_3_lut.init = 16'hcaca;
    LUT4 i24487_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(register_addr[0]), 
         .Z(n30845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24487_3_lut.init = 16'hcaca;
    LUT4 i3847_3_lut (.A(prev_limit_latched), .B(n34347), .C(limit_latched), 
         .Z(n9608)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3847_3_lut.init = 16'hdcdc;
    LUT4 i24665_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i24665_2_lut.init = 16'h9999;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62_adj_373)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[25]), .B(n52), .C(n38), .D(steps_reg[26]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[8]), .B(steps_reg[11]), .C(steps_reg[16]), 
         .D(steps_reg[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(steps_reg[7]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    ClockDivider_U9 step_clk_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .div_factor_reg({div_factor_reg}), .n34347(n34347), .step_clk(step_clk), 
            .n32463(n32463)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (GND_net, debug_c_c, div_factor_reg, n34347, 
            step_clk, n32463) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input n34347;
    output step_clk;
    input n32463;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27328;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n27329, n27327, n32373, n14422, n7160, n7194, n7125;
    wire [31:0]n134;
    
    wire n27674;
    wire [31:0]n40;
    
    wire n27673, n27672, n27671, n27670, n27669, n27668, n27667, 
        n27666, n27665, n27664, n27663, n27662, n27661, n27660, 
        n27659, n27337, n27338, n27336, n27335, n27334, n27333, 
        n27342, n27341, n27332, n27340, n27331, n27330, n27339, 
        n27634, n27633, n27632, n27631, n27630, n27629, n27628, 
        n27627, n27626, n27625, n27624, n27623, n27622, n27621, 
        n27620, n27619, n27614, n27613, n27612, n27611, n27610, 
        n27609, n27608, n27607, n27606, n27605, n27604, n27603, 
        n27602, n27601, n27600, n27599, n27842, n27841, n27840, 
        n27839, n27838, n27837, n27836, n27835, n27834, n27833, 
        n27832, n27831, n27830, n27829, n27828, n27827;
    
    CCU2D sub_1729_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27328), .COUT(n27329));
    defparam sub_1729_add_2_5.INIT0 = 16'h5999;
    defparam sub_1729_add_2_5.INIT1 = 16'h5999;
    defparam sub_1729_add_2_5.INJECT1_0 = "NO";
    defparam sub_1729_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27327), .COUT(n27328));
    defparam sub_1729_add_2_3.INIT0 = 16'h5999;
    defparam sub_1729_add_2_3.INIT1 = 16'h5999;
    defparam sub_1729_add_2_3.INJECT1_0 = "NO";
    defparam sub_1729_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    LUT4 i966_2_lut_rep_248 (.A(n7160), .B(n34347), .Z(n32373)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i966_2_lut_rep_248.init = 16'heeee;
    LUT4 i8656_2_lut_3_lut (.A(n7160), .B(n34347), .C(n7194), .Z(n14422)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8656_2_lut_3_lut.init = 16'he0e0;
    FD1S3IX clk_o_22 (.D(n7125), .CK(debug_c_c), .CD(n32463), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1729_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27327));
    defparam sub_1729_add_2_1.INIT0 = 16'h0000;
    defparam sub_1729_add_2_1.INIT1 = 16'h5999;
    defparam sub_1729_add_2_1.INJECT1_0 = "NO";
    defparam sub_1729_add_2_1.INJECT1_1 = "NO";
    FD1S3IX count_2179__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1S3IX count_2179__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i1.GSR = "ENABLED";
    FD1S3IX count_2179__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i2.GSR = "ENABLED";
    FD1S3IX count_2179__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i3.GSR = "ENABLED";
    FD1S3IX count_2179__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i4.GSR = "ENABLED";
    FD1S3IX count_2179__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i5.GSR = "ENABLED";
    FD1S3IX count_2179__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i6.GSR = "ENABLED";
    FD1S3IX count_2179__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i7.GSR = "ENABLED";
    FD1S3IX count_2179__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i8.GSR = "ENABLED";
    FD1S3IX count_2179__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i9.GSR = "ENABLED";
    FD1S3IX count_2179__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i10.GSR = "ENABLED";
    FD1S3IX count_2179__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i11.GSR = "ENABLED";
    FD1S3IX count_2179__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i12.GSR = "ENABLED";
    FD1S3IX count_2179__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i13.GSR = "ENABLED";
    FD1S3IX count_2179__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i14.GSR = "ENABLED";
    FD1S3IX count_2179__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i15.GSR = "ENABLED";
    FD1S3IX count_2179__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i16.GSR = "ENABLED";
    FD1S3IX count_2179__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i17.GSR = "ENABLED";
    FD1S3IX count_2179__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i18.GSR = "ENABLED";
    FD1S3IX count_2179__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i19.GSR = "ENABLED";
    FD1S3IX count_2179__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i20.GSR = "ENABLED";
    FD1S3IX count_2179__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i21.GSR = "ENABLED";
    FD1S3IX count_2179__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i22.GSR = "ENABLED";
    FD1S3IX count_2179__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i23.GSR = "ENABLED";
    FD1S3IX count_2179__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i24.GSR = "ENABLED";
    FD1S3IX count_2179__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i25.GSR = "ENABLED";
    FD1S3IX count_2179__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i26.GSR = "ENABLED";
    FD1S3IX count_2179__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i27.GSR = "ENABLED";
    FD1S3IX count_2179__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i28.GSR = "ENABLED";
    FD1S3IX count_2179__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i29.GSR = "ENABLED";
    FD1S3IX count_2179__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i30.GSR = "ENABLED";
    FD1S3IX count_2179__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32373), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32373), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32373), .PD(n14422), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27674), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27673), .COUT(n27674), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27672), .COUT(n27673), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27671), .COUT(n27672), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27670), .COUT(n27671), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27669), .COUT(n27670), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27668), .COUT(n27669), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27667), .COUT(n27668), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27666), .COUT(n27667), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27665), .COUT(n27666), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27664), .COUT(n27665), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27663), .COUT(n27664), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27662), .COUT(n27663), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27661), .COUT(n27662), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27660), .COUT(n27661), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27659), .COUT(n27660), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27659), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27337), .COUT(n27338));
    defparam sub_1729_add_2_23.INIT0 = 16'h5999;
    defparam sub_1729_add_2_23.INIT1 = 16'h5999;
    defparam sub_1729_add_2_23.INJECT1_0 = "NO";
    defparam sub_1729_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27336), .COUT(n27337));
    defparam sub_1729_add_2_21.INIT0 = 16'h5999;
    defparam sub_1729_add_2_21.INIT1 = 16'h5999;
    defparam sub_1729_add_2_21.INJECT1_0 = "NO";
    defparam sub_1729_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27335), .COUT(n27336));
    defparam sub_1729_add_2_19.INIT0 = 16'h5999;
    defparam sub_1729_add_2_19.INIT1 = 16'h5999;
    defparam sub_1729_add_2_19.INJECT1_0 = "NO";
    defparam sub_1729_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27334), .COUT(n27335));
    defparam sub_1729_add_2_17.INIT0 = 16'h5999;
    defparam sub_1729_add_2_17.INIT1 = 16'h5999;
    defparam sub_1729_add_2_17.INJECT1_0 = "NO";
    defparam sub_1729_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27333), .COUT(n27334));
    defparam sub_1729_add_2_15.INIT0 = 16'h5999;
    defparam sub_1729_add_2_15.INIT1 = 16'h5999;
    defparam sub_1729_add_2_15.INJECT1_0 = "NO";
    defparam sub_1729_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27342), .S1(n7125));
    defparam sub_1729_add_2_33.INIT0 = 16'h5555;
    defparam sub_1729_add_2_33.INIT1 = 16'h0000;
    defparam sub_1729_add_2_33.INJECT1_0 = "NO";
    defparam sub_1729_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27341), .COUT(n27342));
    defparam sub_1729_add_2_31.INIT0 = 16'h5999;
    defparam sub_1729_add_2_31.INIT1 = 16'h5999;
    defparam sub_1729_add_2_31.INJECT1_0 = "NO";
    defparam sub_1729_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27332), .COUT(n27333));
    defparam sub_1729_add_2_13.INIT0 = 16'h5999;
    defparam sub_1729_add_2_13.INIT1 = 16'h5999;
    defparam sub_1729_add_2_13.INJECT1_0 = "NO";
    defparam sub_1729_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27340), .COUT(n27341));
    defparam sub_1729_add_2_29.INIT0 = 16'h5999;
    defparam sub_1729_add_2_29.INIT1 = 16'h5999;
    defparam sub_1729_add_2_29.INJECT1_0 = "NO";
    defparam sub_1729_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27331), .COUT(n27332));
    defparam sub_1729_add_2_11.INIT0 = 16'h5999;
    defparam sub_1729_add_2_11.INIT1 = 16'h5999;
    defparam sub_1729_add_2_11.INJECT1_0 = "NO";
    defparam sub_1729_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27330), .COUT(n27331));
    defparam sub_1729_add_2_9.INIT0 = 16'h5999;
    defparam sub_1729_add_2_9.INIT1 = 16'h5999;
    defparam sub_1729_add_2_9.INJECT1_0 = "NO";
    defparam sub_1729_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27339), .COUT(n27340));
    defparam sub_1729_add_2_27.INIT0 = 16'h5999;
    defparam sub_1729_add_2_27.INIT1 = 16'h5999;
    defparam sub_1729_add_2_27.INJECT1_0 = "NO";
    defparam sub_1729_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27329), .COUT(n27330));
    defparam sub_1729_add_2_7.INIT0 = 16'h5999;
    defparam sub_1729_add_2_7.INIT1 = 16'h5999;
    defparam sub_1729_add_2_7.INJECT1_0 = "NO";
    defparam sub_1729_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27338), .COUT(n27339));
    defparam sub_1729_add_2_25.INIT0 = 16'h5999;
    defparam sub_1729_add_2_25.INIT1 = 16'h5999;
    defparam sub_1729_add_2_25.INJECT1_0 = "NO";
    defparam sub_1729_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27634), .S1(n7160));
    defparam sub_1731_add_2_33.INIT0 = 16'h5999;
    defparam sub_1731_add_2_33.INIT1 = 16'h0000;
    defparam sub_1731_add_2_33.INJECT1_0 = "NO";
    defparam sub_1731_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27633), .COUT(n27634));
    defparam sub_1731_add_2_31.INIT0 = 16'h5999;
    defparam sub_1731_add_2_31.INIT1 = 16'h5999;
    defparam sub_1731_add_2_31.INJECT1_0 = "NO";
    defparam sub_1731_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27632), .COUT(n27633));
    defparam sub_1731_add_2_29.INIT0 = 16'h5999;
    defparam sub_1731_add_2_29.INIT1 = 16'h5999;
    defparam sub_1731_add_2_29.INJECT1_0 = "NO";
    defparam sub_1731_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27631), .COUT(n27632));
    defparam sub_1731_add_2_27.INIT0 = 16'h5999;
    defparam sub_1731_add_2_27.INIT1 = 16'h5999;
    defparam sub_1731_add_2_27.INJECT1_0 = "NO";
    defparam sub_1731_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27630), .COUT(n27631));
    defparam sub_1731_add_2_25.INIT0 = 16'h5999;
    defparam sub_1731_add_2_25.INIT1 = 16'h5999;
    defparam sub_1731_add_2_25.INJECT1_0 = "NO";
    defparam sub_1731_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27629), .COUT(n27630));
    defparam sub_1731_add_2_23.INIT0 = 16'h5999;
    defparam sub_1731_add_2_23.INIT1 = 16'h5999;
    defparam sub_1731_add_2_23.INJECT1_0 = "NO";
    defparam sub_1731_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27628), .COUT(n27629));
    defparam sub_1731_add_2_21.INIT0 = 16'h5999;
    defparam sub_1731_add_2_21.INIT1 = 16'h5999;
    defparam sub_1731_add_2_21.INJECT1_0 = "NO";
    defparam sub_1731_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27627), .COUT(n27628));
    defparam sub_1731_add_2_19.INIT0 = 16'h5999;
    defparam sub_1731_add_2_19.INIT1 = 16'h5999;
    defparam sub_1731_add_2_19.INJECT1_0 = "NO";
    defparam sub_1731_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27626), .COUT(n27627));
    defparam sub_1731_add_2_17.INIT0 = 16'h5999;
    defparam sub_1731_add_2_17.INIT1 = 16'h5999;
    defparam sub_1731_add_2_17.INJECT1_0 = "NO";
    defparam sub_1731_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27625), .COUT(n27626));
    defparam sub_1731_add_2_15.INIT0 = 16'h5999;
    defparam sub_1731_add_2_15.INIT1 = 16'h5999;
    defparam sub_1731_add_2_15.INJECT1_0 = "NO";
    defparam sub_1731_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27624), .COUT(n27625));
    defparam sub_1731_add_2_13.INIT0 = 16'h5999;
    defparam sub_1731_add_2_13.INIT1 = 16'h5999;
    defparam sub_1731_add_2_13.INJECT1_0 = "NO";
    defparam sub_1731_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27623), .COUT(n27624));
    defparam sub_1731_add_2_11.INIT0 = 16'h5999;
    defparam sub_1731_add_2_11.INIT1 = 16'h5999;
    defparam sub_1731_add_2_11.INJECT1_0 = "NO";
    defparam sub_1731_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27622), .COUT(n27623));
    defparam sub_1731_add_2_9.INIT0 = 16'h5999;
    defparam sub_1731_add_2_9.INIT1 = 16'h5999;
    defparam sub_1731_add_2_9.INJECT1_0 = "NO";
    defparam sub_1731_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27621), .COUT(n27622));
    defparam sub_1731_add_2_7.INIT0 = 16'h5999;
    defparam sub_1731_add_2_7.INIT1 = 16'h5999;
    defparam sub_1731_add_2_7.INJECT1_0 = "NO";
    defparam sub_1731_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27620), .COUT(n27621));
    defparam sub_1731_add_2_5.INIT0 = 16'h5999;
    defparam sub_1731_add_2_5.INIT1 = 16'h5999;
    defparam sub_1731_add_2_5.INJECT1_0 = "NO";
    defparam sub_1731_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27619), .COUT(n27620));
    defparam sub_1731_add_2_3.INIT0 = 16'h5999;
    defparam sub_1731_add_2_3.INIT1 = 16'h5999;
    defparam sub_1731_add_2_3.INJECT1_0 = "NO";
    defparam sub_1731_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27619));
    defparam sub_1731_add_2_1.INIT0 = 16'h0000;
    defparam sub_1731_add_2_1.INIT1 = 16'h5999;
    defparam sub_1731_add_2_1.INJECT1_0 = "NO";
    defparam sub_1731_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27614), .S1(n7194));
    defparam sub_1732_add_2_33.INIT0 = 16'hf555;
    defparam sub_1732_add_2_33.INIT1 = 16'h0000;
    defparam sub_1732_add_2_33.INJECT1_0 = "NO";
    defparam sub_1732_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27613), .COUT(n27614));
    defparam sub_1732_add_2_31.INIT0 = 16'hf555;
    defparam sub_1732_add_2_31.INIT1 = 16'hf555;
    defparam sub_1732_add_2_31.INJECT1_0 = "NO";
    defparam sub_1732_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27612), .COUT(n27613));
    defparam sub_1732_add_2_29.INIT0 = 16'hf555;
    defparam sub_1732_add_2_29.INIT1 = 16'hf555;
    defparam sub_1732_add_2_29.INJECT1_0 = "NO";
    defparam sub_1732_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27611), .COUT(n27612));
    defparam sub_1732_add_2_27.INIT0 = 16'hf555;
    defparam sub_1732_add_2_27.INIT1 = 16'hf555;
    defparam sub_1732_add_2_27.INJECT1_0 = "NO";
    defparam sub_1732_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27610), .COUT(n27611));
    defparam sub_1732_add_2_25.INIT0 = 16'hf555;
    defparam sub_1732_add_2_25.INIT1 = 16'hf555;
    defparam sub_1732_add_2_25.INJECT1_0 = "NO";
    defparam sub_1732_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27609), .COUT(n27610));
    defparam sub_1732_add_2_23.INIT0 = 16'hf555;
    defparam sub_1732_add_2_23.INIT1 = 16'hf555;
    defparam sub_1732_add_2_23.INJECT1_0 = "NO";
    defparam sub_1732_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27608), .COUT(n27609));
    defparam sub_1732_add_2_21.INIT0 = 16'hf555;
    defparam sub_1732_add_2_21.INIT1 = 16'hf555;
    defparam sub_1732_add_2_21.INJECT1_0 = "NO";
    defparam sub_1732_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27607), .COUT(n27608));
    defparam sub_1732_add_2_19.INIT0 = 16'hf555;
    defparam sub_1732_add_2_19.INIT1 = 16'hf555;
    defparam sub_1732_add_2_19.INJECT1_0 = "NO";
    defparam sub_1732_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27606), .COUT(n27607));
    defparam sub_1732_add_2_17.INIT0 = 16'hf555;
    defparam sub_1732_add_2_17.INIT1 = 16'hf555;
    defparam sub_1732_add_2_17.INJECT1_0 = "NO";
    defparam sub_1732_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27605), .COUT(n27606));
    defparam sub_1732_add_2_15.INIT0 = 16'hf555;
    defparam sub_1732_add_2_15.INIT1 = 16'hf555;
    defparam sub_1732_add_2_15.INJECT1_0 = "NO";
    defparam sub_1732_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27604), .COUT(n27605));
    defparam sub_1732_add_2_13.INIT0 = 16'hf555;
    defparam sub_1732_add_2_13.INIT1 = 16'hf555;
    defparam sub_1732_add_2_13.INJECT1_0 = "NO";
    defparam sub_1732_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27603), .COUT(n27604));
    defparam sub_1732_add_2_11.INIT0 = 16'hf555;
    defparam sub_1732_add_2_11.INIT1 = 16'hf555;
    defparam sub_1732_add_2_11.INJECT1_0 = "NO";
    defparam sub_1732_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27602), .COUT(n27603));
    defparam sub_1732_add_2_9.INIT0 = 16'hf555;
    defparam sub_1732_add_2_9.INIT1 = 16'hf555;
    defparam sub_1732_add_2_9.INJECT1_0 = "NO";
    defparam sub_1732_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27601), .COUT(n27602));
    defparam sub_1732_add_2_7.INIT0 = 16'hf555;
    defparam sub_1732_add_2_7.INIT1 = 16'hf555;
    defparam sub_1732_add_2_7.INJECT1_0 = "NO";
    defparam sub_1732_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27600), .COUT(n27601));
    defparam sub_1732_add_2_5.INIT0 = 16'hf555;
    defparam sub_1732_add_2_5.INIT1 = 16'hf555;
    defparam sub_1732_add_2_5.INJECT1_0 = "NO";
    defparam sub_1732_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27599), .COUT(n27600));
    defparam sub_1732_add_2_3.INIT0 = 16'hf555;
    defparam sub_1732_add_2_3.INIT1 = 16'hf555;
    defparam sub_1732_add_2_3.INJECT1_0 = "NO";
    defparam sub_1732_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27599));
    defparam sub_1732_add_2_1.INIT0 = 16'h0000;
    defparam sub_1732_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1732_add_2_1.INJECT1_0 = "NO";
    defparam sub_1732_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27842), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_33.INIT1 = 16'h0000;
    defparam count_2179_add_4_33.INJECT1_0 = "NO";
    defparam count_2179_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27841), .COUT(n27842), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_31.INJECT1_0 = "NO";
    defparam count_2179_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27840), .COUT(n27841), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_29.INJECT1_0 = "NO";
    defparam count_2179_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27839), .COUT(n27840), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_27.INJECT1_0 = "NO";
    defparam count_2179_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27838), .COUT(n27839), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_25.INJECT1_0 = "NO";
    defparam count_2179_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27837), .COUT(n27838), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_23.INJECT1_0 = "NO";
    defparam count_2179_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27836), .COUT(n27837), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_21.INJECT1_0 = "NO";
    defparam count_2179_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27835), .COUT(n27836), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_19.INJECT1_0 = "NO";
    defparam count_2179_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27834), .COUT(n27835), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_17.INJECT1_0 = "NO";
    defparam count_2179_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27833), .COUT(n27834), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_15.INJECT1_0 = "NO";
    defparam count_2179_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27832), .COUT(n27833), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_13.INJECT1_0 = "NO";
    defparam count_2179_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27831), .COUT(n27832), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_11.INJECT1_0 = "NO";
    defparam count_2179_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27830), .COUT(n27831), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_9.INJECT1_0 = "NO";
    defparam count_2179_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27829), .COUT(n27830), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_7.INJECT1_0 = "NO";
    defparam count_2179_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27828), .COUT(n27829), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_5.INJECT1_0 = "NO";
    defparam count_2179_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27827), .COUT(n27828), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_3.INJECT1_0 = "NO";
    defparam count_2179_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27827), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_1.INIT0 = 16'hF000;
    defparam count_2179_add_4_1.INIT1 = 16'h0555;
    defparam count_2179_add_4_1.INJECT1_0 = "NO";
    defparam count_2179_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (\register_addr[1] , databus, 
            n3363, debug_c_c, n34349, VCC_net, GND_net, Stepper_Y_nFault_c, 
            \read_size[0] , Stepper_Y_M0_c_0, n579, \register_addr[0] , 
            n12434, prev_select, n32523, n32509, n32527, n32525, 
            n30283, \select[4] , n32508, n32435, n30454, n32441, 
            n32534, n32449, read_value, n34348, n34351, n34350, 
            n34352, \control_reg[7] , Stepper_Y_En_c, Stepper_Y_Dir_c, 
            Stepper_Y_M2_c_2, Stepper_Y_M1_c_1, \read_size[2] , n30474, 
            n34353, \steps_reg[5] , \steps_reg[3] , n34344, n32420, 
            n34347, n14, n15, limit_c_1, stepping, \register_addr[5] , 
            \register_addr[4] , n32442, rw, n32446, n30450, Stepper_Y_Step_c, 
            n28401, n32463) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[1] ;
    input [31:0]databus;
    input n3363;
    input debug_c_c;
    input n34349;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    output \read_size[0] ;
    output Stepper_Y_M0_c_0;
    input n579;
    input \register_addr[0] ;
    input n12434;
    output prev_select;
    output n32523;
    input n32509;
    input n32527;
    input n32525;
    input n30283;
    input \select[4] ;
    input n32508;
    output n32435;
    input n30454;
    output n32441;
    input n32534;
    output n32449;
    output [31:0]read_value;
    input n34348;
    input n34351;
    input n34350;
    input n34352;
    output \control_reg[7] ;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output Stepper_Y_M2_c_2;
    output Stepper_Y_M1_c_1;
    output \read_size[2] ;
    input n30474;
    input n34353;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input n34344;
    output n32420;
    input n34347;
    input n14;
    input n15;
    input limit_c_1;
    input stepping;
    input \register_addr[5] ;
    input \register_addr[4] ;
    input n32442;
    input rw;
    input n32446;
    input n30450;
    output Stepper_Y_Step_c;
    output n28401;
    input n32463;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30889, n30890, n30891;
    wire [31:0]n224;
    wire [31:0]n3364;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire fault_latched, n12954, n30777, n20514;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n30264, prev_step_clk, step_clk, limit_latched, n182, prev_limit_latched, 
        n32459, n30260, n30275, n30927, n30278, n30270, n32397, 
        n32398, n9612;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n30276, n30883, n30884, int_step, n20526, n32391, n27770, 
        n27769, n27768, n27767, n27766, n27765, n27764, n30925, 
        n27763, n30926, n27762, n18904, n18906, n18907;
    wire [31:0]n5468;
    wire [7:0]n7324;
    wire [31:0]n5432;
    
    wire n27761, n27760, n27759, n27758, n27757, n27756, n5, n6, 
        n27755, n30269, n30258, n49, n41, n60, n54, n42, n62, 
        n52, n38, n58, n50, n56, n46, n30274, n30271, n30277, 
        n30263, n30272, n30257, n30265, n30266, n30267, n30268, 
        n30259, n30256, n30279, n30261, n30262, n30273, n30885;
    
    PFUMX i24533 (.BLUT(n30889), .ALUT(n30890), .C0(\register_addr[1] ), 
          .Z(n30891));
    LUT4 mux_1361_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3363), .Z(n3364[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i1_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i0 (.D(n3364[0]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n30777), .SP(n12954), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n20514), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n30264)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12434), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32459), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i24762_2_lut_3_lut_4_lut_4_lut (.A(n32523), .B(\register_addr[1] ), 
         .C(n32509), .D(n32527), .Z(n30777)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24762_2_lut_3_lut_4_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_365 (.A(div_factor_reg[12]), .B(\register_addr[1] ), 
         .C(steps_reg[12]), .D(\register_addr[0] ), .Z(n30260)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_365.init = 16'hc088;
    LUT4 i13986_3_lut_rep_334_4_lut (.A(n32527), .B(n32525), .C(n30283), 
         .D(\select[4] ), .Z(n32459)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i13986_3_lut_rep_334_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_adj_366 (.A(div_factor_reg[11]), .B(\register_addr[1] ), 
         .C(steps_reg[11]), .D(\register_addr[0] ), .Z(n30275)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_366.init = 16'hc088;
    LUT4 i1_2_lut_rep_310_3_lut_4_lut (.A(n32527), .B(n32525), .C(n32508), 
         .D(\select[4] ), .Z(n32435)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_310_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_316_3_lut_4_lut (.A(n32527), .B(n32525), .C(n30454), 
         .D(\select[4] ), .Z(n32441)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_316_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_324_3_lut_4_lut (.A(n32527), .B(n32525), .C(n32534), 
         .D(\select[4] ), .Z(n32449)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_324_3_lut_4_lut.init = 16'h0100;
    FD1P3IX read_value__i0 (.D(n30927), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_367 (.A(div_factor_reg[10]), .B(\register_addr[1] ), 
         .C(steps_reg[10]), .D(\register_addr[0] ), .Z(n30278)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_367.init = 16'hc088;
    LUT4 i1_4_lut_adj_368 (.A(div_factor_reg[9]), .B(\register_addr[1] ), 
         .C(steps_reg[9]), .D(\register_addr[0] ), .Z(n30270)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_368.init = 16'hc088;
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n32397), .PD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n32397), .PD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n32397), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n32397), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n32397), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n32397), .PD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n32397), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n32397), .PD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n32397), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n32397), .CD(n34350), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n32397), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n32397), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n32398), .CD(n9612), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n32398), .PD(n34352), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n32398), .PD(n34352), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n32398), .CD(n34348), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n32398), .PD(n34352), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n32398), .CD(n34352), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n32398), .PD(n34352), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_369 (.A(div_factor_reg[8]), .B(\register_addr[1] ), 
         .C(steps_reg[8]), .D(\register_addr[0] ), .Z(n30276)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_369.init = 16'hc088;
    FD1P3AX read_size__i2 (.D(n30474), .SP(n12954), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3364[31]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3364[30]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3364[29]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3364[28]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3364[27]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3364[26]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3364[25]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3364[24]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3364[23]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3364[22]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3364[21]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3364[20]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3364[19]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3364[18]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3364[17]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3364[16]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3364[15]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3364[14]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3364[13]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3364[12]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3364[11]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3364[10]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3364[9]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3364[8]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3364[7]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3364[6]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3364[5]), .CK(debug_c_c), .CD(n34353), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3364[4]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3364[3]), .CK(debug_c_c), .CD(n34353), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3364[2]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3364[1]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_295_3_lut (.A(n32459), .B(prev_select), .C(n34344), 
         .Z(n32420)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_295_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n32459), .B(prev_select), .C(n34347), 
         .Z(n12954)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 i24525_3_lut (.A(Stepper_Y_M1_c_1), .B(div_factor_reg[1]), .C(\register_addr[1] ), 
         .Z(n30883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24525_3_lut.init = 16'hcaca;
    LUT4 i24526_3_lut (.A(fault_latched), .B(steps_reg[1]), .C(\register_addr[1] ), 
         .Z(n30884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24526_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n32391), .SP(n20526), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i3851_3_lut (.A(prev_limit_latched), .B(n34347), .C(limit_latched), 
         .Z(n9612)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3851_3_lut.init = 16'hdcdc;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27770), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27769), .COUT(n27770), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27768), .COUT(n27769), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27767), .COUT(n27768), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27766), .COUT(n27767), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27765), .COUT(n27766), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27764), .COUT(n27765), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    LUT4 i24567_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24567_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27763), .COUT(n27764), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    LUT4 i24568_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24568_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27762), .COUT(n27763), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    PFUMX i13166 (.BLUT(n18904), .ALUT(n14), .C0(\register_addr[0] ), 
          .Z(n18906));
    PFUMX i13169 (.BLUT(n18907), .ALUT(n15), .C0(\register_addr[0] ), 
          .Z(n5468[3]));
    LUT4 i14011_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7324[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14011_2_lut.init = 16'h2222;
    LUT4 mux_1620_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5432[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1620_i5_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27761), .COUT(n27762), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27760), .COUT(n27761), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27759), .COUT(n27760), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    LUT4 mux_1361_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3363), 
         .Z(n3364[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i32_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27758), .COUT(n27759), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 i14009_2_lut (.A(\control_reg[7] ), .B(\register_addr[0] ), .Z(n7324[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14009_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27757), .COUT(n27758), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    LUT4 mux_1620_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5432[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1620_i8_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27756), .COUT(n27757), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    PFUMX i6 (.BLUT(n7324[6]), .ALUT(n5), .C0(\register_addr[1] ), .Z(n6));
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27755), .COUT(n27756), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27755), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_1361_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3363), 
         .Z(n3364[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3363), 
         .Z(n3364[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3363), 
         .Z(n3364[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3363), 
         .Z(n3364[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3363), 
         .Z(n3364[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3363), 
         .Z(n3364[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3363), 
         .Z(n3364[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3363), 
         .Z(n3364[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3363), 
         .Z(n3364[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3363), 
         .Z(n3364[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3363), 
         .Z(n3364[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3363), 
         .Z(n3364[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3363), 
         .Z(n3364[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3363), 
         .Z(n3364[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3363), 
         .Z(n3364[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3363), 
         .Z(n3364[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i16_3_lut.init = 16'hcaca;
    LUT4 i24237_2_lut_rep_398 (.A(\register_addr[5] ), .B(\register_addr[4] ), 
         .Z(n32523)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i24237_2_lut_rep_398.init = 16'hbbbb;
    LUT4 i24735_2_lut_4_lut_4_lut (.A(n32442), .B(n34347), .C(n32523), 
         .D(n32420), .Z(n20514)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24735_2_lut_4_lut_4_lut.init = 16'hcdcc;
    LUT4 mux_1361_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3363), 
         .Z(n3364[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3363), 
         .Z(n3364[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3363), 
         .Z(n3364[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3363), 
         .Z(n3364[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3363), 
         .Z(n3364[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3363), .Z(n3364[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3363), .Z(n3364[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3363), .Z(n3364[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3363), .Z(n3364[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3363), .Z(n3364[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3363), .Z(n3364[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3363), .Z(n3364[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3363), .Z(n3364[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3363), .Z(n3364[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_370 (.A(div_factor_reg[22]), .B(\register_addr[1] ), 
         .C(steps_reg[22]), .D(\register_addr[0] ), .Z(n30269)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_370.init = 16'hc088;
    LUT4 i2_3_lut_rep_266 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n32391)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_266.init = 16'h0808;
    LUT4 i14788_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n34347), .Z(n20526)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14788_4_lut_4_lut.init = 16'h0038;
    LUT4 i2_3_lut_rep_272_4_lut (.A(rw), .B(n32446), .C(n30283), .D(n30450), 
         .Z(n32397)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_rep_272_4_lut.init = 16'h4000;
    LUT4 i24742_3_lut_rep_273_3_lut_4_lut (.A(rw), .B(n32446), .C(n32523), 
         .D(n32442), .Z(n32398)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i24742_3_lut_rep_273_3_lut_4_lut.init = 16'h0004;
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12434), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12434), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12434), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12434), .CD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12434), .CD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_371 (.A(div_factor_reg[21]), .B(\register_addr[1] ), 
         .C(steps_reg[21]), .D(\register_addr[0] ), .Z(n30258)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_371.init = 16'hc088;
    LUT4 i17_4_lut (.A(steps_reg[24]), .B(steps_reg[20]), .C(steps_reg[9]), 
         .D(steps_reg[1]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[2]), .B(n52), .C(n38), .D(steps_reg[4]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i26_4_lut.init = 16'hfffe;
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    LUT4 i18_4_lut (.A(steps_reg[0]), .B(steps_reg[10]), .C(steps_reg[28]), 
         .D(\steps_reg[3] ), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[12]), .B(steps_reg[18]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i9_2_lut.init = 16'heeee;
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12434), .CD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12434), .CD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12434), .CD(n34349), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12434), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12434), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12434), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    LUT4 i28_4_lut (.A(steps_reg[22]), .B(n56), .C(n46), .D(\steps_reg[5] ), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_372 (.A(div_factor_reg[20]), .B(\register_addr[1] ), 
         .C(steps_reg[20]), .D(\register_addr[0] ), .Z(n30274)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_372.init = 16'hc088;
    LUT4 i22_4_lut (.A(steps_reg[30]), .B(steps_reg[14]), .C(steps_reg[7]), 
         .D(steps_reg[19]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[16]), .B(steps_reg[27]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i10_2_lut.init = 16'heeee;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12434), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i24_4_lut (.A(steps_reg[23]), .B(steps_reg[13]), .C(steps_reg[29]), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[17]), .B(steps_reg[15]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[21]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[8]), .B(steps_reg[11]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_373 (.A(div_factor_reg[19]), .B(\register_addr[1] ), 
         .C(steps_reg[19]), .D(\register_addr[0] ), .Z(n30271)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_373.init = 16'hc088;
    LUT4 i1_4_lut_adj_374 (.A(div_factor_reg[18]), .B(\register_addr[1] ), 
         .C(steps_reg[18]), .D(\register_addr[0] ), .Z(n30277)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_374.init = 16'hc088;
    LUT4 i13164_3_lut (.A(Stepper_Y_Dir_c), .B(div_factor_reg[5]), .C(\register_addr[1] ), 
         .Z(n18904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13164_3_lut.init = 16'hcaca;
    LUT4 i13167_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(\register_addr[1] ), 
         .Z(n18907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13167_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_375 (.A(div_factor_reg[17]), .B(\register_addr[1] ), 
         .C(steps_reg[17]), .D(\register_addr[0] ), .Z(n30263)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_375.init = 16'hc088;
    LUT4 i1_4_lut_adj_376 (.A(div_factor_reg[16]), .B(\register_addr[1] ), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n30272)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_376.init = 16'hc088;
    FD1P3AX read_value__i31 (.D(n30257), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30265), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30266), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30267), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30268), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n30259), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n30256), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30279), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30264), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30269), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30258), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30274), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30271), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n30277), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n30263), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n30272), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n30261), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30262), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30273), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30260), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n30275), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n30278), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n30270), .SP(n12954), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30276), .SP(n12954), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n5468[7]), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18906), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5468[4]), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5468[3]), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30891), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30885), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i14010_2_lut (.A(Stepper_Y_En_c), .B(\register_addr[0] ), .Z(n7324[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14010_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_377 (.A(div_factor_reg[15]), .B(\register_addr[1] ), 
         .C(steps_reg[15]), .D(\register_addr[0] ), .Z(n30261)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_377.init = 16'hc088;
    LUT4 i1_4_lut_adj_378 (.A(div_factor_reg[14]), .B(\register_addr[1] ), 
         .C(steps_reg[14]), .D(\register_addr[0] ), .Z(n30262)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_378.init = 16'hc088;
    LUT4 i1_4_lut_adj_379 (.A(div_factor_reg[13]), .B(\register_addr[1] ), 
         .C(steps_reg[13]), .D(\register_addr[0] ), .Z(n30273)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_379.init = 16'hc088;
    PFUMX i24527 (.BLUT(n30883), .ALUT(n30884), .C0(\register_addr[0] ), 
          .Z(n30885));
    LUT4 i24671_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i24671_2_lut.init = 16'h9999;
    LUT4 i24531_3_lut (.A(Stepper_Y_M2_c_2), .B(stepping), .C(\register_addr[0] ), 
         .Z(n30889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24531_3_lut.init = 16'hcaca;
    LUT4 i24532_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24532_3_lut.init = 16'hcaca;
    PFUMX i24569 (.BLUT(n30925), .ALUT(n30926), .C0(\register_addr[1] ), 
          .Z(n30927));
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28401)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i31_4_lut.init = 16'hfffe;
    PFUMX mux_1624_i5 (.BLUT(n7324[4]), .ALUT(n5432[4]), .C0(\register_addr[1] ), 
          .Z(n5468[4]));
    PFUMX mux_1624_i8 (.BLUT(n7324[7]), .ALUT(n5432[7]), .C0(\register_addr[1] ), 
          .Z(n5468[7]));
    LUT4 i1_4_lut_adj_380 (.A(div_factor_reg[31]), .B(\register_addr[1] ), 
         .C(steps_reg[31]), .D(\register_addr[0] ), .Z(n30257)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_380.init = 16'hc088;
    LUT4 i1_4_lut_adj_381 (.A(div_factor_reg[30]), .B(\register_addr[1] ), 
         .C(steps_reg[30]), .D(\register_addr[0] ), .Z(n30265)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_381.init = 16'hc088;
    LUT4 i1_4_lut_adj_382 (.A(div_factor_reg[29]), .B(\register_addr[1] ), 
         .C(steps_reg[29]), .D(\register_addr[0] ), .Z(n30266)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_382.init = 16'hc088;
    LUT4 i1_4_lut_adj_383 (.A(div_factor_reg[28]), .B(\register_addr[1] ), 
         .C(steps_reg[28]), .D(\register_addr[0] ), .Z(n30267)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_383.init = 16'hc088;
    LUT4 i1_4_lut_adj_384 (.A(div_factor_reg[27]), .B(\register_addr[1] ), 
         .C(steps_reg[27]), .D(\register_addr[0] ), .Z(n30268)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_384.init = 16'hc088;
    LUT4 i1_4_lut_adj_385 (.A(div_factor_reg[26]), .B(\register_addr[1] ), 
         .C(steps_reg[26]), .D(\register_addr[0] ), .Z(n30259)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_385.init = 16'hc088;
    LUT4 i1_4_lut_adj_386 (.A(div_factor_reg[25]), .B(\register_addr[1] ), 
         .C(steps_reg[25]), .D(\register_addr[0] ), .Z(n30256)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_386.init = 16'hc088;
    LUT4 i1_4_lut_adj_387 (.A(div_factor_reg[24]), .B(\register_addr[1] ), 
         .C(steps_reg[24]), .D(\register_addr[0] ), .Z(n30279)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_387.init = 16'hc088;
    ClockDivider_U7 step_clk_gen (.n34347(n34347), .debug_c_c(debug_c_c), 
            .div_factor_reg({div_factor_reg}), .step_clk(step_clk), .n32463(n32463), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (n34347, debug_c_c, div_factor_reg, step_clk, 
            n32463, GND_net) /* synthesis syn_module_defined=1 */ ;
    input n34347;
    input debug_c_c;
    input [31:0]div_factor_reg;
    output step_clk;
    input n32463;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n6952, n6986, n14396;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n32371, n6917;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27706;
    wire [31:0]n40;
    
    wire n27705, n27704, n27703, n27702, n27701, n27700, n27699, 
        n27698, n27697, n27696, n27695, n27694, n27693, n27692, 
        n27691, n27486, n27485, n27484, n27483, n27482, n27481, 
        n27480, n27479, n27478, n27477, n27476, n27475, n27474, 
        n27473, n27472, n27471, n27470, n27469, n27468, n27467, 
        n27466, n27465, n27464, n27463, n27462, n27461, n27460, 
        n27459, n27458, n27457, n27456, n27455, n27454, n27453, 
        n27452, n27451, n27450, n27449, n27448, n27447, n27446, 
        n27445, n27444, n27443, n27442, n27441, n27440, n27439, 
        n27906, n27905, n27904, n27903, n27902, n27901, n27900, 
        n27899, n27898, n27897, n27896, n27895, n27894, n27893, 
        n27892, n27891;
    
    LUT4 i8630_2_lut_3_lut (.A(n6952), .B(n34347), .C(n6986), .Z(n14396)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8630_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    LUT4 i958_2_lut_rep_246 (.A(n6952), .B(n34347), .Z(n32371)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i958_2_lut_rep_246.init = 16'heeee;
    FD1S3IX clk_o_22 (.D(n6917), .CK(debug_c_c), .CD(n32463), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2177__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i0.GSR = "ENABLED";
    FD1S3IX count_2177__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i1.GSR = "ENABLED";
    FD1S3IX count_2177__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i2.GSR = "ENABLED";
    FD1S3IX count_2177__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i3.GSR = "ENABLED";
    FD1S3IX count_2177__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i4.GSR = "ENABLED";
    FD1S3IX count_2177__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i5.GSR = "ENABLED";
    FD1S3IX count_2177__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i6.GSR = "ENABLED";
    FD1S3IX count_2177__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i7.GSR = "ENABLED";
    FD1S3IX count_2177__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i8.GSR = "ENABLED";
    FD1S3IX count_2177__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i9.GSR = "ENABLED";
    FD1S3IX count_2177__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i10.GSR = "ENABLED";
    FD1S3IX count_2177__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i11.GSR = "ENABLED";
    FD1S3IX count_2177__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i12.GSR = "ENABLED";
    FD1S3IX count_2177__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i13.GSR = "ENABLED";
    FD1S3IX count_2177__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i14.GSR = "ENABLED";
    FD1S3IX count_2177__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i15.GSR = "ENABLED";
    FD1S3IX count_2177__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i16.GSR = "ENABLED";
    FD1S3IX count_2177__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i17.GSR = "ENABLED";
    FD1S3IX count_2177__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i18.GSR = "ENABLED";
    FD1S3IX count_2177__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i19.GSR = "ENABLED";
    FD1S3IX count_2177__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i20.GSR = "ENABLED";
    FD1S3IX count_2177__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i21.GSR = "ENABLED";
    FD1S3IX count_2177__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i22.GSR = "ENABLED";
    FD1S3IX count_2177__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i23.GSR = "ENABLED";
    FD1S3IX count_2177__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i24.GSR = "ENABLED";
    FD1S3IX count_2177__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i25.GSR = "ENABLED";
    FD1S3IX count_2177__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i26.GSR = "ENABLED";
    FD1S3IX count_2177__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i27.GSR = "ENABLED";
    FD1S3IX count_2177__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i28.GSR = "ENABLED";
    FD1S3IX count_2177__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i29.GSR = "ENABLED";
    FD1S3IX count_2177__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i30.GSR = "ENABLED";
    FD1S3IX count_2177__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32371), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i31.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27706), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27705), .COUT(n27706), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27704), .COUT(n27705), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27703), .COUT(n27704), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27702), .COUT(n27703), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27701), .COUT(n27702), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27700), .COUT(n27701), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27699), .COUT(n27700), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27698), .COUT(n27699), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27697), .COUT(n27698), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27696), .COUT(n27697), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27695), .COUT(n27696), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27694), .COUT(n27695), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27693), .COUT(n27694), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27692), .COUT(n27693), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27691), .COUT(n27692), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27691), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    CCU2D sub_1719_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27486), .S1(n6917));
    defparam sub_1719_add_2_33.INIT0 = 16'h5555;
    defparam sub_1719_add_2_33.INIT1 = 16'h0000;
    defparam sub_1719_add_2_33.INJECT1_0 = "NO";
    defparam sub_1719_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27485), .COUT(n27486));
    defparam sub_1719_add_2_31.INIT0 = 16'h5999;
    defparam sub_1719_add_2_31.INIT1 = 16'h5999;
    defparam sub_1719_add_2_31.INJECT1_0 = "NO";
    defparam sub_1719_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    CCU2D sub_1719_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27484), .COUT(n27485));
    defparam sub_1719_add_2_29.INIT0 = 16'h5999;
    defparam sub_1719_add_2_29.INIT1 = 16'h5999;
    defparam sub_1719_add_2_29.INJECT1_0 = "NO";
    defparam sub_1719_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27483), .COUT(n27484));
    defparam sub_1719_add_2_27.INIT0 = 16'h5999;
    defparam sub_1719_add_2_27.INIT1 = 16'h5999;
    defparam sub_1719_add_2_27.INJECT1_0 = "NO";
    defparam sub_1719_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27482), .COUT(n27483));
    defparam sub_1719_add_2_25.INIT0 = 16'h5999;
    defparam sub_1719_add_2_25.INIT1 = 16'h5999;
    defparam sub_1719_add_2_25.INJECT1_0 = "NO";
    defparam sub_1719_add_2_25.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    CCU2D sub_1719_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27481), .COUT(n27482));
    defparam sub_1719_add_2_23.INIT0 = 16'h5999;
    defparam sub_1719_add_2_23.INIT1 = 16'h5999;
    defparam sub_1719_add_2_23.INJECT1_0 = "NO";
    defparam sub_1719_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27480), .COUT(n27481));
    defparam sub_1719_add_2_21.INIT0 = 16'h5999;
    defparam sub_1719_add_2_21.INIT1 = 16'h5999;
    defparam sub_1719_add_2_21.INJECT1_0 = "NO";
    defparam sub_1719_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27479), .COUT(n27480));
    defparam sub_1719_add_2_19.INIT0 = 16'h5999;
    defparam sub_1719_add_2_19.INIT1 = 16'h5999;
    defparam sub_1719_add_2_19.INJECT1_0 = "NO";
    defparam sub_1719_add_2_19.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32371), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    CCU2D sub_1719_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27478), .COUT(n27479));
    defparam sub_1719_add_2_17.INIT0 = 16'h5999;
    defparam sub_1719_add_2_17.INIT1 = 16'h5999;
    defparam sub_1719_add_2_17.INJECT1_0 = "NO";
    defparam sub_1719_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27477), .COUT(n27478));
    defparam sub_1719_add_2_15.INIT0 = 16'h5999;
    defparam sub_1719_add_2_15.INIT1 = 16'h5999;
    defparam sub_1719_add_2_15.INJECT1_0 = "NO";
    defparam sub_1719_add_2_15.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32371), .PD(n14396), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_1719_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27476), .COUT(n27477));
    defparam sub_1719_add_2_13.INIT0 = 16'h5999;
    defparam sub_1719_add_2_13.INIT1 = 16'h5999;
    defparam sub_1719_add_2_13.INJECT1_0 = "NO";
    defparam sub_1719_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27475), .COUT(n27476));
    defparam sub_1719_add_2_11.INIT0 = 16'h5999;
    defparam sub_1719_add_2_11.INIT1 = 16'h5999;
    defparam sub_1719_add_2_11.INJECT1_0 = "NO";
    defparam sub_1719_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27474), .COUT(n27475));
    defparam sub_1719_add_2_9.INIT0 = 16'h5999;
    defparam sub_1719_add_2_9.INIT1 = 16'h5999;
    defparam sub_1719_add_2_9.INJECT1_0 = "NO";
    defparam sub_1719_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27473), .COUT(n27474));
    defparam sub_1719_add_2_7.INIT0 = 16'h5999;
    defparam sub_1719_add_2_7.INIT1 = 16'h5999;
    defparam sub_1719_add_2_7.INJECT1_0 = "NO";
    defparam sub_1719_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27472), .COUT(n27473));
    defparam sub_1719_add_2_5.INIT0 = 16'h5999;
    defparam sub_1719_add_2_5.INIT1 = 16'h5999;
    defparam sub_1719_add_2_5.INJECT1_0 = "NO";
    defparam sub_1719_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27471), .COUT(n27472));
    defparam sub_1719_add_2_3.INIT0 = 16'h5999;
    defparam sub_1719_add_2_3.INIT1 = 16'h5999;
    defparam sub_1719_add_2_3.INJECT1_0 = "NO";
    defparam sub_1719_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27471));
    defparam sub_1719_add_2_1.INIT0 = 16'h0000;
    defparam sub_1719_add_2_1.INIT1 = 16'h5999;
    defparam sub_1719_add_2_1.INJECT1_0 = "NO";
    defparam sub_1719_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27470), .S1(n6952));
    defparam sub_1721_add_2_33.INIT0 = 16'h5999;
    defparam sub_1721_add_2_33.INIT1 = 16'h0000;
    defparam sub_1721_add_2_33.INJECT1_0 = "NO";
    defparam sub_1721_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27469), .COUT(n27470));
    defparam sub_1721_add_2_31.INIT0 = 16'h5999;
    defparam sub_1721_add_2_31.INIT1 = 16'h5999;
    defparam sub_1721_add_2_31.INJECT1_0 = "NO";
    defparam sub_1721_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27468), .COUT(n27469));
    defparam sub_1721_add_2_29.INIT0 = 16'h5999;
    defparam sub_1721_add_2_29.INIT1 = 16'h5999;
    defparam sub_1721_add_2_29.INJECT1_0 = "NO";
    defparam sub_1721_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27467), .COUT(n27468));
    defparam sub_1721_add_2_27.INIT0 = 16'h5999;
    defparam sub_1721_add_2_27.INIT1 = 16'h5999;
    defparam sub_1721_add_2_27.INJECT1_0 = "NO";
    defparam sub_1721_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27466), .COUT(n27467));
    defparam sub_1721_add_2_25.INIT0 = 16'h5999;
    defparam sub_1721_add_2_25.INIT1 = 16'h5999;
    defparam sub_1721_add_2_25.INJECT1_0 = "NO";
    defparam sub_1721_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27465), .COUT(n27466));
    defparam sub_1721_add_2_23.INIT0 = 16'h5999;
    defparam sub_1721_add_2_23.INIT1 = 16'h5999;
    defparam sub_1721_add_2_23.INJECT1_0 = "NO";
    defparam sub_1721_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27464), .COUT(n27465));
    defparam sub_1721_add_2_21.INIT0 = 16'h5999;
    defparam sub_1721_add_2_21.INIT1 = 16'h5999;
    defparam sub_1721_add_2_21.INJECT1_0 = "NO";
    defparam sub_1721_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27463), .COUT(n27464));
    defparam sub_1721_add_2_19.INIT0 = 16'h5999;
    defparam sub_1721_add_2_19.INIT1 = 16'h5999;
    defparam sub_1721_add_2_19.INJECT1_0 = "NO";
    defparam sub_1721_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27462), .COUT(n27463));
    defparam sub_1721_add_2_17.INIT0 = 16'h5999;
    defparam sub_1721_add_2_17.INIT1 = 16'h5999;
    defparam sub_1721_add_2_17.INJECT1_0 = "NO";
    defparam sub_1721_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27461), .COUT(n27462));
    defparam sub_1721_add_2_15.INIT0 = 16'h5999;
    defparam sub_1721_add_2_15.INIT1 = 16'h5999;
    defparam sub_1721_add_2_15.INJECT1_0 = "NO";
    defparam sub_1721_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27460), .COUT(n27461));
    defparam sub_1721_add_2_13.INIT0 = 16'h5999;
    defparam sub_1721_add_2_13.INIT1 = 16'h5999;
    defparam sub_1721_add_2_13.INJECT1_0 = "NO";
    defparam sub_1721_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27459), .COUT(n27460));
    defparam sub_1721_add_2_11.INIT0 = 16'h5999;
    defparam sub_1721_add_2_11.INIT1 = 16'h5999;
    defparam sub_1721_add_2_11.INJECT1_0 = "NO";
    defparam sub_1721_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27458), .COUT(n27459));
    defparam sub_1721_add_2_9.INIT0 = 16'h5999;
    defparam sub_1721_add_2_9.INIT1 = 16'h5999;
    defparam sub_1721_add_2_9.INJECT1_0 = "NO";
    defparam sub_1721_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27457), .COUT(n27458));
    defparam sub_1721_add_2_7.INIT0 = 16'h5999;
    defparam sub_1721_add_2_7.INIT1 = 16'h5999;
    defparam sub_1721_add_2_7.INJECT1_0 = "NO";
    defparam sub_1721_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27456), .COUT(n27457));
    defparam sub_1721_add_2_5.INIT0 = 16'h5999;
    defparam sub_1721_add_2_5.INIT1 = 16'h5999;
    defparam sub_1721_add_2_5.INJECT1_0 = "NO";
    defparam sub_1721_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27455), .COUT(n27456));
    defparam sub_1721_add_2_3.INIT0 = 16'h5999;
    defparam sub_1721_add_2_3.INIT1 = 16'h5999;
    defparam sub_1721_add_2_3.INJECT1_0 = "NO";
    defparam sub_1721_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27455));
    defparam sub_1721_add_2_1.INIT0 = 16'h0000;
    defparam sub_1721_add_2_1.INIT1 = 16'h5999;
    defparam sub_1721_add_2_1.INJECT1_0 = "NO";
    defparam sub_1721_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27454), .S1(n6986));
    defparam sub_1722_add_2_33.INIT0 = 16'hf555;
    defparam sub_1722_add_2_33.INIT1 = 16'h0000;
    defparam sub_1722_add_2_33.INJECT1_0 = "NO";
    defparam sub_1722_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27453), .COUT(n27454));
    defparam sub_1722_add_2_31.INIT0 = 16'hf555;
    defparam sub_1722_add_2_31.INIT1 = 16'hf555;
    defparam sub_1722_add_2_31.INJECT1_0 = "NO";
    defparam sub_1722_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27452), .COUT(n27453));
    defparam sub_1722_add_2_29.INIT0 = 16'hf555;
    defparam sub_1722_add_2_29.INIT1 = 16'hf555;
    defparam sub_1722_add_2_29.INJECT1_0 = "NO";
    defparam sub_1722_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27451), .COUT(n27452));
    defparam sub_1722_add_2_27.INIT0 = 16'hf555;
    defparam sub_1722_add_2_27.INIT1 = 16'hf555;
    defparam sub_1722_add_2_27.INJECT1_0 = "NO";
    defparam sub_1722_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27450), .COUT(n27451));
    defparam sub_1722_add_2_25.INIT0 = 16'hf555;
    defparam sub_1722_add_2_25.INIT1 = 16'hf555;
    defparam sub_1722_add_2_25.INJECT1_0 = "NO";
    defparam sub_1722_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27449), .COUT(n27450));
    defparam sub_1722_add_2_23.INIT0 = 16'hf555;
    defparam sub_1722_add_2_23.INIT1 = 16'hf555;
    defparam sub_1722_add_2_23.INJECT1_0 = "NO";
    defparam sub_1722_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27448), .COUT(n27449));
    defparam sub_1722_add_2_21.INIT0 = 16'hf555;
    defparam sub_1722_add_2_21.INIT1 = 16'hf555;
    defparam sub_1722_add_2_21.INJECT1_0 = "NO";
    defparam sub_1722_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27447), .COUT(n27448));
    defparam sub_1722_add_2_19.INIT0 = 16'hf555;
    defparam sub_1722_add_2_19.INIT1 = 16'hf555;
    defparam sub_1722_add_2_19.INJECT1_0 = "NO";
    defparam sub_1722_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27446), .COUT(n27447));
    defparam sub_1722_add_2_17.INIT0 = 16'hf555;
    defparam sub_1722_add_2_17.INIT1 = 16'hf555;
    defparam sub_1722_add_2_17.INJECT1_0 = "NO";
    defparam sub_1722_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27445), .COUT(n27446));
    defparam sub_1722_add_2_15.INIT0 = 16'hf555;
    defparam sub_1722_add_2_15.INIT1 = 16'hf555;
    defparam sub_1722_add_2_15.INJECT1_0 = "NO";
    defparam sub_1722_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27444), .COUT(n27445));
    defparam sub_1722_add_2_13.INIT0 = 16'hf555;
    defparam sub_1722_add_2_13.INIT1 = 16'hf555;
    defparam sub_1722_add_2_13.INJECT1_0 = "NO";
    defparam sub_1722_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27443), .COUT(n27444));
    defparam sub_1722_add_2_11.INIT0 = 16'hf555;
    defparam sub_1722_add_2_11.INIT1 = 16'hf555;
    defparam sub_1722_add_2_11.INJECT1_0 = "NO";
    defparam sub_1722_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27442), .COUT(n27443));
    defparam sub_1722_add_2_9.INIT0 = 16'hf555;
    defparam sub_1722_add_2_9.INIT1 = 16'hf555;
    defparam sub_1722_add_2_9.INJECT1_0 = "NO";
    defparam sub_1722_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27441), .COUT(n27442));
    defparam sub_1722_add_2_7.INIT0 = 16'hf555;
    defparam sub_1722_add_2_7.INIT1 = 16'hf555;
    defparam sub_1722_add_2_7.INJECT1_0 = "NO";
    defparam sub_1722_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27440), .COUT(n27441));
    defparam sub_1722_add_2_5.INIT0 = 16'hf555;
    defparam sub_1722_add_2_5.INIT1 = 16'hf555;
    defparam sub_1722_add_2_5.INJECT1_0 = "NO";
    defparam sub_1722_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27439), .COUT(n27440));
    defparam sub_1722_add_2_3.INIT0 = 16'hf555;
    defparam sub_1722_add_2_3.INIT1 = 16'hf555;
    defparam sub_1722_add_2_3.INJECT1_0 = "NO";
    defparam sub_1722_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27439));
    defparam sub_1722_add_2_1.INIT0 = 16'h0000;
    defparam sub_1722_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1722_add_2_1.INJECT1_0 = "NO";
    defparam sub_1722_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27906), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_33.INIT1 = 16'h0000;
    defparam count_2177_add_4_33.INJECT1_0 = "NO";
    defparam count_2177_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27905), .COUT(n27906), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_31.INJECT1_0 = "NO";
    defparam count_2177_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27904), .COUT(n27905), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_29.INJECT1_0 = "NO";
    defparam count_2177_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27903), .COUT(n27904), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_27.INJECT1_0 = "NO";
    defparam count_2177_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27902), .COUT(n27903), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_25.INJECT1_0 = "NO";
    defparam count_2177_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27901), .COUT(n27902), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_23.INJECT1_0 = "NO";
    defparam count_2177_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27900), .COUT(n27901), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_21.INJECT1_0 = "NO";
    defparam count_2177_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27899), .COUT(n27900), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_19.INJECT1_0 = "NO";
    defparam count_2177_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27898), .COUT(n27899), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_17.INJECT1_0 = "NO";
    defparam count_2177_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27897), .COUT(n27898), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_15.INJECT1_0 = "NO";
    defparam count_2177_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27896), .COUT(n27897), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_13.INJECT1_0 = "NO";
    defparam count_2177_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27895), .COUT(n27896), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_11.INJECT1_0 = "NO";
    defparam count_2177_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27894), .COUT(n27895), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_9.INJECT1_0 = "NO";
    defparam count_2177_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27893), .COUT(n27894), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_7.INJECT1_0 = "NO";
    defparam count_2177_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27892), .COUT(n27893), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_5.INJECT1_0 = "NO";
    defparam count_2177_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27891), .COUT(n27892), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_3.INJECT1_0 = "NO";
    defparam count_2177_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27891), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_1.INIT0 = 16'hF000;
    defparam count_2177_add_4_1.INIT1 = 16'h0555;
    defparam count_2177_add_4_1.INJECT1_0 = "NO";
    defparam count_2177_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (\register_addr[0] , databus_out, n2, rw, databus, 
            \read_value[13] , n1, n32503, \read_value[13]_adj_43 , read_value, 
            n32407, n52, n2_adj_45, \read_value[12]_adj_46 , n1_adj_47, 
            \read_value[12]_adj_48 , \register_addr[2] , \register_addr[1] , 
            n2_adj_49, \select[7] , n32527, n32509, n30454, n30363, 
            n32523, n30474, n32534, n30658, n29690, n30435, n2_adj_50, 
            \read_value[11]_adj_51 , n1_adj_52, \read_value[11]_adj_53 , 
            n2_adj_54, \read_value[10]_adj_55 , n1_adj_56, \read_value[10]_adj_57 , 
            \register_addr[4] , n2_adj_58, \read_value[18]_adj_59 , n1_adj_60, 
            \read_value[18]_adj_61 , \read_size[0] , \read_size[0]_adj_62 , 
            \register_addr[5] , \read_size[0]_adj_63 , \read_size[0]_adj_64 , 
            read_size, \select[1] , n32511, \sendcount[1] , n11271, 
            n2_adj_66, \read_value[19]_adj_67 , n1_adj_68, \read_value[9]_adj_69 , 
            n1_adj_70, n2_adj_71, \read_value[25]_adj_72 , n1_adj_73, 
            n2_adj_74, \read_value[9]_adj_75 , \read_value[19]_adj_76 , 
            n2_adj_77, \read_value[17]_adj_78 , n1_adj_79, \read_value[17]_adj_80 , 
            n2_adj_81, \read_value[20]_adj_82 , n1_adj_83, \read_value[16]_adj_84 , 
            n1_adj_85, \read_value[16]_adj_86 , \read_value[25]_adj_87 , 
            n32486, \register_addr[3] , n30594, n2_adj_88, \read_value[15]_adj_89 , 
            n1_adj_90, n2_adj_91, \read_value[15]_adj_92 , \read_value[8]_adj_93 , 
            n1_adj_94, n2_adj_95, \read_value[14]_adj_96 , n1_adj_97, 
            n2_adj_98, \read_value[14]_adj_99 , \read_value[30]_adj_100 , 
            n1_adj_101, n32416, n30450, n32379, \read_value[8]_adj_102 , 
            n2_adj_103, \select[2] , \read_size[0]_adj_104 , n5, n32469, 
            n6, \reg_size[2] , \read_value[24]_adj_105 , n1_adj_106, 
            \read_value[24]_adj_107 , \read_value[20]_adj_108 , n4, \read_value[7]_adj_109 , 
            n32406, \read_value[7]_adj_110 , \read_value[7]_adj_111 , 
            n32408, n34344, read_value_adj_186, n64, n4_adj_120, \read_value[6]_adj_121 , 
            \read_value[6]_adj_122 , \read_value[6]_adj_123 , \read_value[30]_adj_124 , 
            n2_adj_125, \read_value[23]_adj_126 , n1_adj_127, n4_adj_128, 
            \read_value[23]_adj_129 , \read_value[5]_adj_130 , \read_value[5]_adj_131 , 
            \read_value[5]_adj_132 , n4_adj_133, \read_value[4]_adj_134 , 
            \read_value[4]_adj_135 , \read_value[4]_adj_136 , n2_adj_137, 
            \read_value[22]_adj_138 , n1_adj_139, n2_adj_140, \read_value[29]_adj_141 , 
            n1_adj_142, \read_value[22]_adj_143 , \read_size[2]_adj_144 , 
            \read_size[2]_adj_145 , \read_size[2]_adj_146 , \read_size[2]_adj_147 , 
            n4_adj_148, \read_value[3]_adj_149 , \read_value[3]_adj_150 , 
            \read_value[3]_adj_151 , n2_adj_152, \read_value[31]_adj_153 , 
            n1_adj_154, \read_value[31]_adj_155 , n2_adj_156, n4_adj_157, 
            \read_value[2]_adj_158 , \read_value[2]_adj_159 , \read_value[2]_adj_160 , 
            \read_value[28]_adj_161 , n1_adj_162, \read_value[28]_adj_163 , 
            n1_adj_164, \read_value[1]_adj_165 , n6_adj_166, \read_value[1]_adj_167 , 
            n4_adj_168, \read_value[0]_adj_169 , \read_value[0]_adj_170 , 
            \read_value[0]_adj_171 , \read_value[29]_adj_172 , n2_adj_173, 
            n2_adj_174, \read_value[27]_adj_175 , n1_adj_176, \read_value[21]_adj_177 , 
            n1_adj_178, \read_value[27]_adj_179 , n2_adj_180, \read_value[26]_adj_181 , 
            n1_adj_182, \read_value[26]_adj_183 , \read_value[21]_adj_184 , 
            n31057, debug_c_c, n28352, GND_net, n32375, rc_ch8_c, 
            n12030, n30942, n28337, n31041, rc_ch7_c, n12031, n31025, 
            n11987, n34347, n31050, rc_ch4_c, n30958, n28331, n12138, 
            n28345, n30999, rc_ch3_c, n31033, n32369, n14446, n1000, 
            n988, rc_ch2_c, n54, n4_adj_185, n32374, n31079, n28339, 
            rc_ch1_c, n30940) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[0] ;
    input [31:0]databus_out;
    input n2;
    input rw;
    output [31:0]databus;
    input \read_value[13] ;
    input n1;
    input n32503;
    input \read_value[13]_adj_43 ;
    input [31:0]read_value;
    input n32407;
    input n52;
    input n2_adj_45;
    input \read_value[12]_adj_46 ;
    input n1_adj_47;
    input \read_value[12]_adj_48 ;
    input \register_addr[2] ;
    input \register_addr[1] ;
    input n2_adj_49;
    input \select[7] ;
    input n32527;
    input n32509;
    output n30454;
    output n30363;
    input n32523;
    output n30474;
    output n32534;
    output n30658;
    output n29690;
    output n30435;
    input n2_adj_50;
    input \read_value[11]_adj_51 ;
    input n1_adj_52;
    input \read_value[11]_adj_53 ;
    input n2_adj_54;
    input \read_value[10]_adj_55 ;
    input n1_adj_56;
    input \read_value[10]_adj_57 ;
    input \register_addr[4] ;
    input n2_adj_58;
    input \read_value[18]_adj_59 ;
    input n1_adj_60;
    input \read_value[18]_adj_61 ;
    input \read_size[0] ;
    input \read_size[0]_adj_62 ;
    input \register_addr[5] ;
    input \read_size[0]_adj_63 ;
    input \read_size[0]_adj_64 ;
    input [2:0]read_size;
    input \select[1] ;
    output n32511;
    input \sendcount[1] ;
    output n11271;
    input n2_adj_66;
    input \read_value[19]_adj_67 ;
    input n1_adj_68;
    input \read_value[9]_adj_69 ;
    input n1_adj_70;
    input n2_adj_71;
    input \read_value[25]_adj_72 ;
    input n1_adj_73;
    input n2_adj_74;
    input \read_value[9]_adj_75 ;
    input \read_value[19]_adj_76 ;
    input n2_adj_77;
    input \read_value[17]_adj_78 ;
    input n1_adj_79;
    input \read_value[17]_adj_80 ;
    input n2_adj_81;
    input \read_value[20]_adj_82 ;
    input n1_adj_83;
    input \read_value[16]_adj_84 ;
    input n1_adj_85;
    input \read_value[16]_adj_86 ;
    input \read_value[25]_adj_87 ;
    input n32486;
    input \register_addr[3] ;
    input n30594;
    input n2_adj_88;
    input \read_value[15]_adj_89 ;
    input n1_adj_90;
    input n2_adj_91;
    input \read_value[15]_adj_92 ;
    input \read_value[8]_adj_93 ;
    input n1_adj_94;
    input n2_adj_95;
    input \read_value[14]_adj_96 ;
    input n1_adj_97;
    input n2_adj_98;
    input \read_value[14]_adj_99 ;
    input \read_value[30]_adj_100 ;
    input n1_adj_101;
    input n32416;
    input n30450;
    output n32379;
    input \read_value[8]_adj_102 ;
    input n2_adj_103;
    input \select[2] ;
    input \read_size[0]_adj_104 ;
    output n5;
    input n32469;
    output n6;
    output \reg_size[2] ;
    input \read_value[24]_adj_105 ;
    input n1_adj_106;
    input \read_value[24]_adj_107 ;
    input \read_value[20]_adj_108 ;
    input n4;
    input \read_value[7]_adj_109 ;
    input n32406;
    input \read_value[7]_adj_110 ;
    input \read_value[7]_adj_111 ;
    input n32408;
    input n34344;
    input [7:0]read_value_adj_186;
    input n64;
    input n4_adj_120;
    input \read_value[6]_adj_121 ;
    input \read_value[6]_adj_122 ;
    input \read_value[6]_adj_123 ;
    input \read_value[30]_adj_124 ;
    input n2_adj_125;
    input \read_value[23]_adj_126 ;
    input n1_adj_127;
    input n4_adj_128;
    input \read_value[23]_adj_129 ;
    input \read_value[5]_adj_130 ;
    input \read_value[5]_adj_131 ;
    input \read_value[5]_adj_132 ;
    input n4_adj_133;
    input \read_value[4]_adj_134 ;
    input \read_value[4]_adj_135 ;
    input \read_value[4]_adj_136 ;
    input n2_adj_137;
    input \read_value[22]_adj_138 ;
    input n1_adj_139;
    input n2_adj_140;
    input \read_value[29]_adj_141 ;
    input n1_adj_142;
    input \read_value[22]_adj_143 ;
    input \read_size[2]_adj_144 ;
    input \read_size[2]_adj_145 ;
    input \read_size[2]_adj_146 ;
    input \read_size[2]_adj_147 ;
    input n4_adj_148;
    input \read_value[3]_adj_149 ;
    input \read_value[3]_adj_150 ;
    input \read_value[3]_adj_151 ;
    input n2_adj_152;
    input \read_value[31]_adj_153 ;
    input n1_adj_154;
    input \read_value[31]_adj_155 ;
    input n2_adj_156;
    input n4_adj_157;
    input \read_value[2]_adj_158 ;
    input \read_value[2]_adj_159 ;
    input \read_value[2]_adj_160 ;
    input \read_value[28]_adj_161 ;
    input n1_adj_162;
    input \read_value[28]_adj_163 ;
    input n1_adj_164;
    input \read_value[1]_adj_165 ;
    input n6_adj_166;
    input \read_value[1]_adj_167 ;
    input n4_adj_168;
    input \read_value[0]_adj_169 ;
    input \read_value[0]_adj_170 ;
    input \read_value[0]_adj_171 ;
    input \read_value[29]_adj_172 ;
    input n2_adj_173;
    input n2_adj_174;
    input \read_value[27]_adj_175 ;
    input n1_adj_176;
    input \read_value[21]_adj_177 ;
    input n1_adj_178;
    input \read_value[27]_adj_179 ;
    input n2_adj_180;
    input \read_value[26]_adj_181 ;
    input n1_adj_182;
    input \read_value[26]_adj_183 ;
    input \read_value[21]_adj_184 ;
    output n31057;
    input debug_c_c;
    input n28352;
    input GND_net;
    input n32375;
    input rc_ch8_c;
    input n12030;
    output n30942;
    input n28337;
    output n31041;
    input rc_ch7_c;
    input n12031;
    output n31025;
    input n11987;
    input n34347;
    output n31050;
    input rc_ch4_c;
    output n30958;
    input n28331;
    input n12138;
    input n28345;
    output n30999;
    input rc_ch3_c;
    output n31033;
    input n32369;
    input n14446;
    output n1000;
    output n988;
    input rc_ch2_c;
    output n54;
    output n4_adj_185;
    input n32374;
    output n31079;
    input n28339;
    input rc_ch1_c;
    output n30940;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n979;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n31529, n1039, n32231, n10, n8;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n32227;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n32228, n10_adj_137, n32266, n8_adj_139, n32267, n31807, 
        n31804, n31808;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n32269, n31806, n31805, n1009, n32270, n10_adj_143, n32284, 
        n31803, n31802, n32283, n32286, n32287;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(213[12:21])
    
    wire n176, n10_adj_145, n8_adj_147, n31526, n31525, n31527, 
        n10_adj_151, n8_adj_153, n19, n22, n25, n32314, n32313, 
        n32316, n31774, n31771, n31775, n32317, n10_adj_157, n8_adj_159, 
        n31773, n31772, n31528, n32504;
    wire [7:0]read_value_adj_368;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(212[12:22])
    
    wire n7, n7_adj_163, n7_adj_164, n7_adj_165, n7_adj_166, n7_adj_167, 
        n7_adj_168, n32354, n18, n21, n24, n32353, n32356, n994, 
        n32357, n31770, n31769, n10_adj_173, n8_adj_175, n8_adj_177, 
        n10_adj_179, n8_adj_181, n10_adj_183, n10_adj_189, n8_adj_191, 
        n10_adj_195, n8_adj_197, n8_adj_199, n32460, n31531, n10_adj_205, 
        n8_adj_207, n10_adj_209, n8_adj_213, n10_adj_215, n8_adj_217, 
        n10_adj_219, n8_adj_223, n32230, n32233, n32319, n32289, 
        n32272, n32359, n10_adj_227, n8_adj_231, n32358, n32355, 
        n13, n12, n6_adj_237, n10_adj_239, n13_adj_244, n12_adj_246, 
        n6_adj_247, n10_adj_249, n10_adj_256, n32318, n32315, n8_adj_258, 
        n13_adj_260, n12_adj_262, n6_adj_263, n10_adj_267, n13_adj_270, 
        n12_adj_272, n6_adj_273, n10_adj_275, n10_adj_282, n8_adj_284, 
        n10_adj_286, n32288, n32285, n8_adj_288, n13_adj_296, n12_adj_298, 
        n6_adj_299, n10_adj_301, n10_adj_304, n8_adj_308, n1024, n10_adj_312, 
        n13_adj_314, n12_adj_316, n6_adj_317, n10_adj_319, n32271, 
        n32268, n8_adj_322, n14, n10_adj_329, n7_adj_330, n12_adj_332, 
        n32232, n32229, n13_adj_337, n12_adj_339, n6_adj_340, n10_adj_342, 
        n10_adj_349, n10_adj_351, n8_adj_353, n31530, n8_adj_355, 
        n10_adj_359, n8_adj_361, n1054;
    
    LUT4 n979_bdd_3_lut_25225 (.A(n979), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n31529)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n979_bdd_3_lut_25225.init = 16'he2e2;
    LUT4 n1039_bdd_3_lut_25198 (.A(n1039), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n32231)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1039_bdd_3_lut_25198.init = 16'he2e2;
    LUT4 i5_4_lut (.A(databus_out[13]), .B(n10), .C(n2), .D(rw), .Z(databus[13])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfcfe;
    LUT4 i4_4_lut (.A(\read_value[13] ), .B(n8), .C(n1), .D(n32503), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_25202 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n32227)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25202.init = 16'h2222;
    LUT4 i2_4_lut (.A(\read_value[13]_adj_43 ), .B(read_value[13]), .C(n32407), 
         .D(n52), .Z(n8)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_25203 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n32228)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25203.init = 16'he4e4;
    LUT4 i5_4_lut_adj_261 (.A(databus_out[12]), .B(n10_adj_137), .C(n2_adj_45), 
         .D(rw), .Z(databus[12])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_261.init = 16'hfcfe;
    LUT4 register_addr_1__bdd_2_lut_25213 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n32266)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25213.init = 16'h2222;
    LUT4 i4_4_lut_adj_262 (.A(\read_value[12]_adj_46 ), .B(n8_adj_139), 
         .C(n1_adj_47), .D(n32503), .Z(n10_adj_137)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_262.init = 16'hfefc;
    LUT4 i2_4_lut_adj_263 (.A(\read_value[12]_adj_48 ), .B(read_value[12]), 
         .C(n32407), .D(n52), .Z(n8_adj_139)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_263.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_25214 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n32267)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25214.init = 16'he4e4;
    L6MUX21 i25056 (.D0(n31807), .D1(n31804), .SD(\register_addr[2] ), 
            .Z(n31808));
    LUT4 n1009_bdd_3_lut_25208 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n32269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1009_bdd_3_lut_25208.init = 16'hcaca;
    PFUMX i25054 (.BLUT(n31806), .ALUT(n31805), .C0(\register_addr[1] ), 
          .Z(n31807));
    LUT4 n1009_bdd_3_lut_26007 (.A(n1009), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n32270)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1009_bdd_3_lut_26007.init = 16'he2e2;
    LUT4 i5_4_lut_adj_264 (.A(databus_out[19]), .B(n10_adj_143), .C(n2_adj_49), 
         .D(rw), .Z(databus[19])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_264.init = 16'hfcfe;
    LUT4 register_addr_1__bdd_3_lut_25233 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n32284)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25233.init = 16'he4e4;
    PFUMX i25051 (.BLUT(n31803), .ALUT(n31802), .C0(\register_addr[1] ), 
          .Z(n31804));
    LUT4 register_addr_1__bdd_2_lut_25232 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n32283)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25232.init = 16'h2222;
    LUT4 \register_1[[4__bdd_3_lut_25984  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n32286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_25984 .init = 16'hcaca;
    LUT4 \register_1[[4__bdd_2_lut_25985  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n32287)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_25985 .init = 16'h8888;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32527), .B(n32509), .C(n30454), .D(\register_addr[1] ), 
         .Z(n30363)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_265 (.A(n32527), .B(n32509), .C(n32523), 
         .D(\register_addr[1] ), .Z(n30474)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_265.init = 16'h0100;
    LUT4 i24836_2_lut_3_lut_4_lut (.A(n32527), .B(n32509), .C(\register_addr[1] ), 
         .D(n32534), .Z(n30658)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24836_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_266 (.A(n32527), .B(n32509), .C(\register_addr[1] ), 
         .D(n32534), .Z(n29690)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_266.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_267 (.A(n32527), .B(n32509), .C(n30454), 
         .D(\register_addr[1] ), .Z(n30435)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_267.init = 16'h0010;
    LUT4 i5_4_lut_adj_268 (.A(databus_out[11]), .B(n10_adj_145), .C(n2_adj_50), 
         .D(rw), .Z(databus[11])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_268.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_269 (.A(\read_value[11]_adj_51 ), .B(n8_adj_147), 
         .C(n1_adj_52), .D(n32503), .Z(n10_adj_145)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_269.init = 16'hfefc;
    PFUMX i24940 (.BLUT(n31526), .ALUT(n31525), .C0(\register_addr[1] ), 
          .Z(n31527));
    LUT4 i2_4_lut_adj_270 (.A(\read_value[11]_adj_53 ), .B(read_value[11]), 
         .C(n32407), .D(n52), .Z(n8_adj_147)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_270.init = 16'heca0;
    LUT4 i5_4_lut_adj_271 (.A(databus_out[10]), .B(n10_adj_151), .C(n2_adj_54), 
         .D(rw), .Z(databus[10])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_271.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_272 (.A(\read_value[10]_adj_55 ), .B(n8_adj_153), 
         .C(n1_adj_56), .D(n32503), .Z(n10_adj_151)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_272.init = 16'hfefc;
    LUT4 i2_4_lut_adj_273 (.A(\read_value[10]_adj_57 ), .B(read_value[10]), 
         .C(n32407), .D(n52), .Z(n8_adj_153)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_273.init = 16'heca0;
    PFUMX i38 (.BLUT(n19), .ALUT(n22), .C0(\register_addr[4] ), .Z(n25));
    LUT4 register_addr_1__bdd_3_lut_25264 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n32314)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25264.init = 16'he4e4;
    LUT4 register_addr_1__bdd_3_lut_25023 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n31526)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25023.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_25263 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n32313)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25263.init = 16'h2222;
    LUT4 \register_1[[5__bdd_3_lut_25908  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n32316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_25908 .init = 16'hcaca;
    L6MUX21 i25031 (.D0(n31774), .D1(n31771), .SD(\register_addr[2] ), 
            .Z(n31775));
    LUT4 \register_1[[5__bdd_2_lut_25909  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n32317)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_25909 .init = 16'h8888;
    LUT4 register_addr_1__bdd_2_lut_25022 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n31525)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25022.init = 16'h2222;
    LUT4 i5_4_lut_adj_274 (.A(databus_out[18]), .B(n10_adj_157), .C(n2_adj_58), 
         .D(rw), .Z(databus[18])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_274.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_275 (.A(\read_value[18]_adj_59 ), .B(n8_adj_159), 
         .C(n1_adj_60), .D(n32503), .Z(n10_adj_157)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_275.init = 16'hfefc;
    LUT4 i2_4_lut_adj_276 (.A(\read_value[18]_adj_61 ), .B(read_value[18]), 
         .C(n32407), .D(n52), .Z(n8_adj_159)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_276.init = 16'heca0;
    PFUMX i25029 (.BLUT(n31773), .ALUT(n31772), .C0(\register_addr[1] ), 
          .Z(n31774));
    LUT4 n979_bdd_3_lut_24942 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n31528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n979_bdd_3_lut_24942.init = 16'hcaca;
    LUT4 i14_2_lut_rep_379 (.A(\select[7] ), .B(rw), .Z(n32504)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam i14_2_lut_rep_379.init = 16'h8888;
    LUT4 Select_3620_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[5]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3620_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3619_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[6]), 
         .Z(n7_adj_163)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3619_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3618_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[7]), 
         .Z(n7_adj_164)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3618_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3625_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[0]), 
         .Z(n7_adj_165)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3625_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3623_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[2]), 
         .Z(n7_adj_166)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3623_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3622_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[3]), 
         .Z(n7_adj_167)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3622_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3621_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[4]), 
         .Z(n7_adj_168)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3621_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 i24570_3_lut (.A(\read_size[0] ), .B(\read_size[0]_adj_62 ), .C(\register_addr[5] ), 
         .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24570_3_lut.init = 16'hcaca;
    LUT4 i24571_3_lut (.A(\read_size[0]_adj_63 ), .B(\read_size[0]_adj_64 ), 
         .C(\register_addr[5] ), .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24571_3_lut.init = 16'hcaca;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n32354)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    PFUMX i37 (.BLUT(n18), .ALUT(n21), .C0(\register_addr[4] ), .Z(n24));
    LUT4 Select_3633_i1_2_lut_rep_386 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n32511)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3633_i1_2_lut_rep_386.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n11271)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n32353)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    LUT4 n994_bdd_3_lut_25272 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n32356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n994_bdd_3_lut_25272.init = 16'hcaca;
    LUT4 n994_bdd_3_lut_25882 (.A(n994), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n32357)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n994_bdd_3_lut_25882.init = 16'he2e2;
    PFUMX i25026 (.BLUT(n31770), .ALUT(n31769), .C0(\register_addr[1] ), 
          .Z(n31771));
    LUT4 i5_4_lut_adj_277 (.A(databus_out[9]), .B(n10_adj_173), .C(n2_adj_66), 
         .D(rw), .Z(databus[9])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_277.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_278 (.A(\read_value[19]_adj_67 ), .B(n8_adj_175), 
         .C(n1_adj_68), .D(n32503), .Z(n10_adj_143)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_278.init = 16'hfefc;
    LUT4 i4_4_lut_adj_279 (.A(\read_value[9]_adj_69 ), .B(n8_adj_177), .C(n1_adj_70), 
         .D(n32503), .Z(n10_adj_173)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_279.init = 16'hfefc;
    LUT4 i5_4_lut_adj_280 (.A(databus_out[25]), .B(n10_adj_179), .C(n2_adj_71), 
         .D(rw), .Z(databus[25])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_280.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_281 (.A(\read_value[25]_adj_72 ), .B(n8_adj_181), 
         .C(n1_adj_73), .D(n32503), .Z(n10_adj_179)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_281.init = 16'hfefc;
    LUT4 i5_4_lut_adj_282 (.A(databus_out[20]), .B(n10_adj_183), .C(n2_adj_74), 
         .D(rw), .Z(databus[20])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_282.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_283 (.A(\read_value[9]_adj_75 ), .B(read_value[9]), 
         .C(n32407), .D(n52), .Z(n8_adj_177)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_283.init = 16'heca0;
    LUT4 i2_4_lut_adj_284 (.A(\read_value[19]_adj_76 ), .B(read_value[19]), 
         .C(n32407), .D(n52), .Z(n8_adj_175)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_284.init = 16'heca0;
    LUT4 i5_4_lut_adj_285 (.A(databus_out[17]), .B(n10_adj_189), .C(n2_adj_77), 
         .D(rw), .Z(databus[17])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_285.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_286 (.A(\read_value[17]_adj_78 ), .B(n8_adj_191), 
         .C(n1_adj_79), .D(n32503), .Z(n10_adj_189)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_286.init = 16'hfefc;
    LUT4 i2_4_lut_adj_287 (.A(\read_value[17]_adj_80 ), .B(read_value[17]), 
         .C(n32407), .D(n52), .Z(n8_adj_191)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_287.init = 16'heca0;
    LUT4 i5_4_lut_adj_288 (.A(databus_out[16]), .B(n10_adj_195), .C(n2_adj_81), 
         .D(rw), .Z(databus[16])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_288.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_289 (.A(\read_value[20]_adj_82 ), .B(n8_adj_197), 
         .C(n1_adj_83), .D(n32503), .Z(n10_adj_183)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_289.init = 16'hfefc;
    LUT4 i4_4_lut_adj_290 (.A(\read_value[16]_adj_84 ), .B(n8_adj_199), 
         .C(n1_adj_85), .D(n32503), .Z(n10_adj_195)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_290.init = 16'hfefc;
    LUT4 i2_4_lut_adj_291 (.A(\read_value[16]_adj_86 ), .B(read_value[16]), 
         .C(n32407), .D(n52), .Z(n8_adj_199)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_291.init = 16'heca0;
    FD1S3IX read_value__i0 (.D(n31531), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_292 (.A(\read_value[25]_adj_87 ), .B(read_value[25]), 
         .C(n32407), .D(n52), .Z(n8_adj_181)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_292.init = 16'heca0;
    LUT4 i2_4_lut_rep_335 (.A(n32486), .B(\register_addr[2] ), .C(\register_addr[3] ), 
         .D(n30594), .Z(n32460)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(221[7:31])
    defparam i2_4_lut_rep_335.init = 16'hfefa;
    LUT4 i14584_1_lut_4_lut (.A(n32486), .B(\register_addr[2] ), .C(\register_addr[3] ), 
         .D(n30594), .Z(n176)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(221[7:31])
    defparam i14584_1_lut_4_lut.init = 16'h0105;
    LUT4 i5_4_lut_adj_293 (.A(databus_out[15]), .B(n10_adj_205), .C(n2_adj_88), 
         .D(rw), .Z(databus[15])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_293.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_294 (.A(\read_value[15]_adj_89 ), .B(n8_adj_207), 
         .C(n1_adj_90), .D(n32503), .Z(n10_adj_205)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_294.init = 16'hfefc;
    LUT4 i5_4_lut_adj_295 (.A(databus_out[8]), .B(n10_adj_209), .C(n2_adj_91), 
         .D(rw), .Z(databus[8])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_295.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_296 (.A(\read_value[15]_adj_92 ), .B(read_value[15]), 
         .C(n32407), .D(n52), .Z(n8_adj_207)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_296.init = 16'heca0;
    LUT4 i4_4_lut_adj_297 (.A(\read_value[8]_adj_93 ), .B(n8_adj_213), .C(n1_adj_94), 
         .D(n32503), .Z(n10_adj_209)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_297.init = 16'hfefc;
    LUT4 i24246_2_lut_rep_409 (.A(\register_addr[4] ), .B(\register_addr[5] ), 
         .Z(n32534)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i24246_2_lut_rep_409.init = 16'hbbbb;
    LUT4 i5_4_lut_adj_298 (.A(databus_out[14]), .B(n10_adj_215), .C(n2_adj_95), 
         .D(rw), .Z(databus[14])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_298.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_299 (.A(\read_value[14]_adj_96 ), .B(n8_adj_217), 
         .C(n1_adj_97), .D(n32503), .Z(n10_adj_215)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_299.init = 16'hfefc;
    LUT4 i5_4_lut_adj_300 (.A(databus_out[30]), .B(n10_adj_219), .C(n2_adj_98), 
         .D(rw), .Z(databus[30])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_300.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_301 (.A(\read_value[14]_adj_99 ), .B(read_value[14]), 
         .C(n32407), .D(n52), .Z(n8_adj_217)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_301.init = 16'heca0;
    LUT4 i4_4_lut_adj_302 (.A(\read_value[30]_adj_100 ), .B(n8_adj_223), 
         .C(n1_adj_101), .D(n32503), .Z(n10_adj_219)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_302.init = 16'hfefc;
    LUT4 i1_2_lut_rep_254_4_lut (.A(rw), .B(n30454), .C(n32416), .D(n30450), 
         .Z(n32379)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_254_4_lut.init = 16'h4000;
    LUT4 n1039_bdd_3_lut_25190 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n32230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1039_bdd_3_lut_25190.init = 16'hcaca;
    LUT4 i2_4_lut_adj_303 (.A(\read_value[8]_adj_102 ), .B(read_value[8]), 
         .C(n32407), .D(n52), .Z(n8_adj_213)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_303.init = 16'heca0;
    FD1S3IX read_value__i7 (.D(n31808), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\register_addr[4] ), .B(\register_addr[5] ), .Z(n30454)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    FD1S3IX read_value__i6 (.D(n32233), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n32319), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n32289), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n31775), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n32272), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i1 (.D(n32359), .CK(\select[7] ), .CD(n32460), 
            .Q(read_value_adj_368[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_304 (.A(databus_out[24]), .B(n10_adj_227), .C(n2_adj_103), 
         .D(rw), .Z(databus[24])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_304.init = 16'hfcfe;
    LUT4 i1_4_lut (.A(\select[2] ), .B(read_size_c[0]), .C(\read_size[0]_adj_104 ), 
         .D(\select[7] ), .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i2_4_lut_adj_305 (.A(read_size[0]), .B(n25), .C(\select[1] ), 
         .D(n32469), .Z(n6)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_305.init = 16'heca0;
    LUT4 i1_4_lut_adj_306 (.A(read_size[2]), .B(n24), .C(\select[1] ), 
         .D(n32469), .Z(\reg_size[2] )) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_306.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_25040 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n31770)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25040.init = 16'he4e4;
    LUT4 i4_4_lut_adj_307 (.A(\read_value[24]_adj_105 ), .B(n8_adj_231), 
         .C(n1_adj_106), .D(n32503), .Z(n10_adj_227)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_307.init = 16'hfefc;
    LUT4 i2_4_lut_adj_308 (.A(\read_value[24]_adj_107 ), .B(read_value[24]), 
         .C(n32407), .D(n52), .Z(n8_adj_231)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_308.init = 16'heca0;
    LUT4 i2_4_lut_adj_309 (.A(\read_value[20]_adj_108 ), .B(read_value[20]), 
         .C(n32407), .D(n52), .Z(n8_adj_197)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_309.init = 16'heca0;
    L6MUX21 i25275 (.D0(n32358), .D1(n32355), .SD(\register_addr[2] ), 
            .Z(n32359));
    PFUMX i25273 (.BLUT(n32357), .ALUT(n32356), .C0(\register_addr[1] ), 
          .Z(n32358));
    PFUMX i25270 (.BLUT(n32354), .ALUT(n32353), .C0(\register_addr[1] ), 
          .Z(n32355));
    LUT4 i7_4_lut (.A(n13), .B(n4), .C(n12), .D(n6_adj_237), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut_adj_310 (.A(\read_value[7]_adj_109 ), .B(n10_adj_239), 
         .C(n7_adj_164), .D(n32406), .Z(n13)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_310.init = 16'hfefc;
    LUT4 i4_4_lut_adj_311 (.A(\read_value[7]_adj_110 ), .B(\read_value[7]_adj_111 ), 
         .C(n32408), .D(n32503), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_311.init = 16'heca0;
    LUT4 Select_3618_i6_2_lut (.A(databus_out[7]), .B(n34344), .Z(n6_adj_237)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3618_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_312 (.A(read_value[7]), .B(read_value_adj_186[7]), 
         .C(n52), .D(n64), .Z(n10_adj_239)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_312.init = 16'heca0;
    LUT4 i7_4_lut_adj_313 (.A(n13_adj_244), .B(n4_adj_120), .C(n12_adj_246), 
         .D(n6_adj_247), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_313.init = 16'hfffe;
    LUT4 i5_4_lut_adj_314 (.A(\read_value[6]_adj_121 ), .B(n10_adj_249), 
         .C(n7_adj_163), .D(n32406), .Z(n13_adj_244)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_314.init = 16'hfefc;
    LUT4 i4_4_lut_adj_315 (.A(\read_value[6]_adj_122 ), .B(\read_value[6]_adj_123 ), 
         .C(n32408), .D(n32503), .Z(n12_adj_246)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_315.init = 16'heca0;
    LUT4 Select_3619_i6_2_lut (.A(databus_out[6]), .B(n34344), .Z(n6_adj_247)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3619_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_316 (.A(read_value[6]), .B(read_value_adj_186[6]), 
         .C(n52), .D(n64), .Z(n10_adj_249)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_316.init = 16'heca0;
    LUT4 i2_4_lut_adj_317 (.A(\read_value[30]_adj_124 ), .B(read_value[30]), 
         .C(n32407), .D(n52), .Z(n8_adj_223)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_317.init = 16'heca0;
    LUT4 i5_4_lut_adj_318 (.A(databus_out[23]), .B(n10_adj_256), .C(n2_adj_125), 
         .D(rw), .Z(databus[23])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_318.init = 16'hfcfe;
    L6MUX21 i25242 (.D0(n32318), .D1(n32315), .SD(\register_addr[2] ), 
            .Z(n32319));
    LUT4 i4_4_lut_adj_319 (.A(\read_value[23]_adj_126 ), .B(n8_adj_258), 
         .C(n1_adj_127), .D(n32503), .Z(n10_adj_256)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_319.init = 16'hfefc;
    PFUMX i25240 (.BLUT(n32317), .ALUT(n32316), .C0(\register_addr[1] ), 
          .Z(n32318));
    LUT4 i7_4_lut_adj_320 (.A(n13_adj_260), .B(n4_adj_128), .C(n12_adj_262), 
         .D(n6_adj_263), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_320.init = 16'hfffe;
    PFUMX i25238 (.BLUT(n32314), .ALUT(n32313), .C0(\register_addr[1] ), 
          .Z(n32315));
    LUT4 i2_4_lut_adj_321 (.A(\read_value[23]_adj_129 ), .B(read_value[23]), 
         .C(n32407), .D(n52), .Z(n8_adj_258)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_321.init = 16'heca0;
    LUT4 i5_4_lut_adj_322 (.A(\read_value[5]_adj_130 ), .B(n10_adj_267), 
         .C(n7), .D(n32406), .Z(n13_adj_260)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_322.init = 16'hfefc;
    LUT4 i4_4_lut_adj_323 (.A(\read_value[5]_adj_131 ), .B(\read_value[5]_adj_132 ), 
         .C(n32408), .D(n32503), .Z(n12_adj_262)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_323.init = 16'heca0;
    LUT4 i7_4_lut_adj_324 (.A(n13_adj_270), .B(n4_adj_133), .C(n12_adj_272), 
         .D(n6_adj_273), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_324.init = 16'hfffe;
    LUT4 Select_3620_i6_2_lut (.A(databus_out[5]), .B(rw), .Z(n6_adj_263)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3620_i6_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_325 (.A(\read_value[4]_adj_134 ), .B(n10_adj_275), 
         .C(n7_adj_168), .D(n32406), .Z(n13_adj_270)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_325.init = 16'hfefc;
    LUT4 i2_4_lut_adj_326 (.A(read_value[5]), .B(read_value_adj_186[5]), 
         .C(n52), .D(n64), .Z(n10_adj_267)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_326.init = 16'heca0;
    LUT4 i4_4_lut_adj_327 (.A(\read_value[4]_adj_135 ), .B(\read_value[4]_adj_136 ), 
         .C(n32408), .D(n32503), .Z(n12_adj_272)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_327.init = 16'heca0;
    LUT4 Select_3621_i6_2_lut (.A(databus_out[4]), .B(rw), .Z(n6_adj_273)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3621_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_328 (.A(read_value[4]), .B(read_value_adj_186[4]), 
         .C(n52), .D(n64), .Z(n10_adj_275)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_328.init = 16'heca0;
    LUT4 i5_4_lut_adj_329 (.A(databus_out[22]), .B(n10_adj_282), .C(n2_adj_137), 
         .D(rw), .Z(databus[22])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_329.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_330 (.A(\read_value[22]_adj_138 ), .B(n8_adj_284), 
         .C(n1_adj_139), .D(n32503), .Z(n10_adj_282)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_330.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_25039 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n31769)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25039.init = 16'h2222;
    LUT4 i5_4_lut_adj_331 (.A(databus_out[29]), .B(n10_adj_286), .C(n2_adj_140), 
         .D(rw), .Z(databus[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_331.init = 16'hfcfe;
    L6MUX21 i25221 (.D0(n32288), .D1(n32285), .SD(\register_addr[2] ), 
            .Z(n32289));
    LUT4 i4_4_lut_adj_332 (.A(\read_value[29]_adj_141 ), .B(n8_adj_288), 
         .C(n1_adj_142), .D(n32503), .Z(n10_adj_286)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_332.init = 16'hfefc;
    LUT4 i2_4_lut_adj_333 (.A(\read_value[22]_adj_143 ), .B(read_value[22]), 
         .C(n32407), .D(n52), .Z(n8_adj_284)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_333.init = 16'heca0;
    LUT4 i39_3_lut (.A(\read_size[2]_adj_144 ), .B(\read_size[2]_adj_145 ), 
         .C(\register_addr[5] ), .Z(n18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i39_3_lut.init = 16'hcaca;
    LUT4 i38_3_lut (.A(\read_size[2]_adj_146 ), .B(\read_size[2]_adj_147 ), 
         .C(\register_addr[5] ), .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38_3_lut.init = 16'hcaca;
    LUT4 i7_4_lut_adj_334 (.A(n13_adj_296), .B(n4_adj_148), .C(n12_adj_298), 
         .D(n6_adj_299), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_334.init = 16'hfffe;
    PFUMX i25219 (.BLUT(n32287), .ALUT(n32286), .C0(\register_addr[1] ), 
          .Z(n32288));
    LUT4 i5_4_lut_adj_335 (.A(\read_value[3]_adj_149 ), .B(n10_adj_301), 
         .C(n7_adj_167), .D(n32406), .Z(n13_adj_296)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_335.init = 16'hfefc;
    LUT4 i4_4_lut_adj_336 (.A(\read_value[3]_adj_150 ), .B(\read_value[3]_adj_151 ), 
         .C(n32408), .D(n32503), .Z(n12_adj_298)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_336.init = 16'heca0;
    PFUMX i25217 (.BLUT(n32284), .ALUT(n32283), .C0(\register_addr[1] ), 
          .Z(n32285));
    LUT4 Select_3622_i6_2_lut (.A(databus_out[3]), .B(rw), .Z(n6_adj_299)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3622_i6_2_lut.init = 16'h2222;
    LUT4 n1024_bdd_3_lut_25028 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n31772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1024_bdd_3_lut_25028.init = 16'hcaca;
    LUT4 i5_4_lut_adj_337 (.A(databus_out[31]), .B(n10_adj_304), .C(n2_adj_152), 
         .D(rw), .Z(databus[31])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_337.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_338 (.A(read_value[3]), .B(read_value_adj_186[3]), 
         .C(n52), .D(n64), .Z(n10_adj_301)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_338.init = 16'heca0;
    LUT4 i4_4_lut_adj_339 (.A(\read_value[31]_adj_153 ), .B(n8_adj_308), 
         .C(n1_adj_154), .D(n32503), .Z(n10_adj_304)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_339.init = 16'hfefc;
    LUT4 i2_4_lut_adj_340 (.A(\read_value[31]_adj_155 ), .B(read_value[31]), 
         .C(n32407), .D(n52), .Z(n8_adj_308)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_340.init = 16'heca0;
    LUT4 n1024_bdd_3_lut_25639 (.A(n1024), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n31773)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1024_bdd_3_lut_25639.init = 16'he2e2;
    LUT4 i5_4_lut_adj_341 (.A(databus_out[28]), .B(n10_adj_312), .C(n2_adj_156), 
         .D(rw), .Z(databus[28])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_341.init = 16'hfcfe;
    LUT4 i7_4_lut_adj_342 (.A(n13_adj_314), .B(n4_adj_157), .C(n12_adj_316), 
         .D(n6_adj_317), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_342.init = 16'hfffe;
    LUT4 i5_4_lut_adj_343 (.A(\read_value[2]_adj_158 ), .B(n10_adj_319), 
         .C(n7_adj_166), .D(n32406), .Z(n13_adj_314)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_343.init = 16'hfefc;
    LUT4 i4_4_lut_adj_344 (.A(\read_value[2]_adj_159 ), .B(\read_value[2]_adj_160 ), 
         .C(n32408), .D(n32503), .Z(n12_adj_316)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_344.init = 16'heca0;
    L6MUX21 i25211 (.D0(n32271), .D1(n32268), .SD(\register_addr[2] ), 
            .Z(n32272));
    LUT4 i4_4_lut_adj_345 (.A(\read_value[28]_adj_161 ), .B(n8_adj_322), 
         .C(n1_adj_162), .D(n32503), .Z(n10_adj_312)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_345.init = 16'hfefc;
    LUT4 Select_3623_i6_2_lut (.A(databus_out[2]), .B(rw), .Z(n6_adj_317)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3623_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_346 (.A(read_value[2]), .B(read_value_adj_186[2]), 
         .C(n52), .D(n64), .Z(n10_adj_319)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_346.init = 16'heca0;
    PFUMX i25209 (.BLUT(n32270), .ALUT(n32269), .C0(\register_addr[1] ), 
          .Z(n32271));
    LUT4 i2_4_lut_adj_347 (.A(\read_value[28]_adj_163 ), .B(read_value[28]), 
         .C(n32407), .D(n52), .Z(n8_adj_322)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_347.init = 16'heca0;
    PFUMX i25206 (.BLUT(n32267), .ALUT(n32266), .C0(\register_addr[1] ), 
          .Z(n32268));
    LUT4 i7_4_lut_adj_348 (.A(n1_adj_164), .B(n14), .C(n10_adj_329), .D(n7_adj_330), 
         .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_348.init = 16'hfffe;
    LUT4 i6_4_lut (.A(\read_value[1]_adj_165 ), .B(n12_adj_332), .C(n6_adj_166), 
         .D(n32407), .Z(n14)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    L6MUX21 i25193 (.D0(n32232), .D1(n32229), .SD(\register_addr[2] ), 
            .Z(n32233));
    LUT4 i2_4_lut_adj_349 (.A(read_value[1]), .B(read_value_adj_186[1]), 
         .C(n52), .D(n64), .Z(n10_adj_329)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_349.init = 16'heca0;
    LUT4 Select_3624_i7_2_lut (.A(databus_out[1]), .B(rw), .Z(n7_adj_330)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3624_i7_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_350 (.A(\read_value[1]_adj_167 ), .B(read_value_adj_368[1]), 
         .C(n32408), .D(n32504), .Z(n12_adj_332)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_350.init = 16'heca0;
    PFUMX i25191 (.BLUT(n32231), .ALUT(n32230), .C0(\register_addr[1] ), 
          .Z(n32232));
    LUT4 i7_4_lut_adj_351 (.A(n13_adj_337), .B(n4_adj_168), .C(n12_adj_339), 
         .D(n6_adj_340), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_351.init = 16'hfffe;
    LUT4 i5_4_lut_adj_352 (.A(\read_value[0]_adj_169 ), .B(n10_adj_342), 
         .C(n7_adj_165), .D(n32406), .Z(n13_adj_337)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_352.init = 16'hfefc;
    LUT4 i4_4_lut_adj_353 (.A(\read_value[0]_adj_170 ), .B(\read_value[0]_adj_171 ), 
         .C(n32408), .D(n32503), .Z(n12_adj_339)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_353.init = 16'heca0;
    LUT4 Select_3625_i6_2_lut (.A(databus_out[0]), .B(n34344), .Z(n6_adj_340)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3625_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_354 (.A(read_value[0]), .B(read_value_adj_186[0]), 
         .C(n52), .D(n64), .Z(n10_adj_342)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_354.init = 16'heca0;
    PFUMX i25188 (.BLUT(n32228), .ALUT(n32227), .C0(\register_addr[1] ), 
          .Z(n32229));
    LUT4 i2_4_lut_adj_355 (.A(\read_value[29]_adj_172 ), .B(read_value[29]), 
         .C(n32407), .D(n52), .Z(n8_adj_288)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_355.init = 16'heca0;
    LUT4 i5_4_lut_adj_356 (.A(databus_out[21]), .B(n10_adj_349), .C(n2_adj_173), 
         .D(rw), .Z(databus[21])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_356.init = 16'hfcfe;
    LUT4 i5_4_lut_adj_357 (.A(databus_out[27]), .B(n10_adj_351), .C(n2_adj_174), 
         .D(rw), .Z(databus[27])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_357.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_358 (.A(\read_value[27]_adj_175 ), .B(n8_adj_353), 
         .C(n1_adj_176), .D(n32503), .Z(n10_adj_351)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_358.init = 16'hfefc;
    L6MUX21 i24945 (.D0(n31530), .D1(n31527), .SD(\register_addr[2] ), 
            .Z(n31531));
    LUT4 i4_4_lut_adj_359 (.A(\read_value[21]_adj_177 ), .B(n8_adj_355), 
         .C(n1_adj_178), .D(n32503), .Z(n10_adj_349)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_359.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_25129 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n31803)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25129.init = 16'he4e4;
    LUT4 i2_4_lut_adj_360 (.A(\read_value[27]_adj_179 ), .B(read_value[27]), 
         .C(n32407), .D(n52), .Z(n8_adj_353)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_360.init = 16'heca0;
    LUT4 i5_4_lut_adj_361 (.A(databus_out[26]), .B(n10_adj_359), .C(n2_adj_180), 
         .D(rw), .Z(databus[26])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_361.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_362 (.A(\read_value[26]_adj_181 ), .B(n8_adj_361), 
         .C(n1_adj_182), .D(n32503), .Z(n10_adj_359)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_362.init = 16'hfefc;
    LUT4 i2_4_lut_adj_363 (.A(\read_value[26]_adj_183 ), .B(read_value[26]), 
         .C(n32407), .D(n52), .Z(n8_adj_361)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_363.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_25128 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n31802)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25128.init = 16'h2222;
    PFUMX i24943 (.BLUT(n31529), .ALUT(n31528), .C0(\register_addr[1] ), 
          .Z(n31530));
    LUT4 i2_4_lut_adj_364 (.A(\read_value[21]_adj_184 ), .B(read_value[21]), 
         .C(n32407), .D(n52), .Z(n8_adj_355)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_364.init = 16'heca0;
    LUT4 n1054_bdd_3_lut_25053 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n31805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1054_bdd_3_lut_25053.init = 16'hcaca;
    LUT4 n1054_bdd_3_lut_25375 (.A(n1054), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n31806)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1054_bdd_3_lut_25375.init = 16'he2e2;
    PWMReceiver recv_ch8 (.n31057(n31057), .n1054(n1054), .debug_c_c(debug_c_c), 
            .n28352(n28352), .GND_net(GND_net), .n32375(n32375), .rc_ch8_c(rc_ch8_c), 
            .\register[6] ({\register[6] }), .n12030(n12030), .n30942(n30942)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(259[14] 263[36])
    PWMReceiver_U1 recv_ch7 (.n1039(n1039), .debug_c_c(debug_c_c), .n28337(n28337), 
            .GND_net(GND_net), .n31041(n31041), .n32375(n32375), .rc_ch7_c(rc_ch7_c), 
            .\register[5] ({\register[5] }), .n12031(n12031), .n31025(n31025)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(254[14] 258[36])
    PWMReceiver_U2 recv_ch4 (.\register[4] ({\register[4] }), .debug_c_c(debug_c_c), 
            .n11987(n11987), .n32375(n32375), .GND_net(GND_net), .n34347(n34347), 
            .n31050(n31050), .rc_ch4_c(rc_ch4_c), .n30958(n30958), .n1024(n1024), 
            .n28331(n28331)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(249[14] 253[36])
    PWMReceiver_U3 recv_ch3 (.debug_c_c(debug_c_c), .n32375(n32375), .GND_net(GND_net), 
            .\register[3] ({\register[3] }), .n12138(n12138), .n1009(n1009), 
            .n28345(n28345), .n30999(n30999), .rc_ch3_c(rc_ch3_c), .n31033(n31033)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(244[14] 248[36])
    PWMReceiver_U4 recv_ch2 (.debug_c_c(debug_c_c), .n32375(n32375), .GND_net(GND_net), 
            .\register[2] ({\register[2] }), .n32369(n32369), .n14446(n14446), 
            .n994(n994), .n1000(n1000), .n988(n988), .rc_ch2_c(rc_ch2_c), 
            .n54(n54), .n4(n4_adj_185)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(239[14] 243[36])
    PWMReceiver_U5 recv_ch1 (.debug_c_c(debug_c_c), .n32375(n32375), .GND_net(GND_net), 
            .\register[1] ({\register[1] }), .n32374(n32374), .n31079(n31079), 
            .n979(n979), .n28339(n28339), .rc_ch1_c(rc_ch1_c), .n30940(n30940)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(234[17] 238[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (n31057, n1054, debug_c_c, n28352, GND_net, n32375, 
            rc_ch8_c, \register[6] , n12030, n30942) /* synthesis syn_module_defined=1 */ ;
    output n31057;
    output n1054;
    input debug_c_c;
    input n28352;
    input GND_net;
    input n32375;
    input rc_ch8_c;
    output [7:0]\register[6] ;
    input n12030;
    output n30942;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n32487, n11840, n32419, n30461, n28200, n10, n30679, 
        n32421, n30507, n32399, n30525, n32533, n32526, n28430, 
        n28349, n32524, n30175, n54, n32448, n30140, n32470, n4, 
        n32530, n1048, n1060, n20263, n28382, n32529, n6, n30526, 
        n32528, n32485, n4_adj_133, n32483, n4_adj_134, n32484, 
        n28511;
    wire [7:0]n943;
    wire [7:0]n43;
    
    wire n32447, n30737;
    wire [15:0]n116;
    
    wire n14198, n27350, n27349, n27348, n27347, n27346, n27345, 
        n27344, n27343, n27638, n27637, n27636, n27635, n12;
    
    LUT4 i1_2_lut_rep_294_3_lut_4_lut (.A(count[12]), .B(n32487), .C(count[9]), 
         .D(n11840), .Z(n32419)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_294_3_lut_4_lut.init = 16'hfffe;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n32419), .C(n30461), 
         .D(n28200), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i24323_3_lut_4_lut (.A(count[8]), .B(n32419), .C(n28200), .D(n30461), 
         .Z(n30679)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i24323_3_lut_4_lut.init = 16'hfeee;
    LUT4 i24805_3_lut_4_lut_4_lut (.A(n32421), .B(n30507), .C(n32399), 
         .D(n28200), .Z(n30525)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i24805_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i24790_4_lut (.A(n32533), .B(n32526), .C(n28430), .D(n28349), 
         .Z(n31057)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i24790_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n30679), .B(n32524), .C(n11840), .D(n30175), .Z(n28349)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 i3_4_lut (.A(n54), .B(n32448), .C(n30140), .D(n32470), .Z(n30175)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n11840)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(count[4]), .B(count[5]), .C(n4), .D(n32530), .Z(n28200)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut.init = 16'hc800;
    LUT4 i5_2_lut_rep_401 (.A(n1048), .B(n1060), .Z(n32526)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_401.init = 16'h4444;
    LUT4 i3_4_lut_adj_255 (.A(count[7]), .B(count[8]), .C(n20263), .D(count[6]), 
         .Z(n28382)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_255.init = 16'hfffe;
    LUT4 i14534_4_lut (.A(count[0]), .B(n32529), .C(n6), .D(count[3]), 
         .Z(n20263)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i14534_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1048), .B(n1060), .C(n28430), .D(n32533), 
         .Z(n30526)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_4_lut_adj_256 (.A(n32419), .B(count[8]), .C(n32528), .D(n32485), 
         .Z(n30140)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_256.init = 16'hfbbb;
    LUT4 i2_4_lut_adj_257 (.A(count[13]), .B(count[12]), .C(n11840), .D(n4_adj_133), 
         .Z(n28430)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_257.init = 16'h8880;
    LUT4 i1_4_lut_adj_258 (.A(count[5]), .B(count[9]), .C(n32483), .D(n4_adj_134), 
         .Z(n4_adj_133)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_258.init = 16'hfcec;
    LUT4 i3_3_lut_4_lut (.A(count[8]), .B(n32530), .C(n32484), .D(n32529), 
         .Z(n28511)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_259 (.A(n32529), .B(n32530), .C(n32528), 
         .D(count[0]), .Z(n30461)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_259.init = 16'h8000;
    LUT4 i14268_2_lut (.A(n943[0]), .B(n30140), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14268_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_322_3_lut_4_lut (.A(n32533), .B(count[13]), .C(n11840), 
         .D(count[12]), .Z(n32447)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_322_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX valid_48 (.D(n30525), .SP(n28352), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1054));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_274_3_lut_4_lut (.A(n11840), .B(n32470), .C(count[8]), 
         .D(count[9]), .Z(n32399)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_274_3_lut_4_lut.init = 16'hfffe;
    LUT4 i14754_2_lut_rep_323 (.A(n28382), .B(count[9]), .Z(n32448)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14754_2_lut_rep_323.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_260 (.A(n28382), .B(count[9]), .C(n32470), 
         .D(n11840), .Z(n30507)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_260.init = 16'hfff8;
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n32375), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1060));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1060), .SP(n32375), .CK(debug_c_c), .Q(n1048));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_399 (.A(n1060), .B(n1048), .Z(n32524)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_399.init = 16'hbbbb;
    LUT4 i24379_2_lut_3_lut_4_lut (.A(n1060), .B(n1048), .C(count[13]), 
         .D(n32533), .Z(n30737)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i24379_2_lut_3_lut_4_lut.init = 16'hfffb;
    LUT4 i2_3_lut_rep_403 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n32528)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_403.init = 16'h8080;
    LUT4 i1_2_lut_rep_359_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n32484)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_359_4_lut.init = 16'h8000;
    LUT4 i14050_2_lut_rep_404 (.A(count[5]), .B(count[4]), .Z(n32529)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14050_2_lut_rep_404.init = 16'h8888;
    LUT4 i1_2_lut_rep_405 (.A(count[6]), .B(count[7]), .Z(n32530)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_405.init = 16'h8888;
    LUT4 i1_2_lut_rep_358_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n32483)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_358_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_rep_360_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[4]), 
         .D(count[5]), .Z(n32485)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_rep_360_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_134)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_408 (.A(count[15]), .B(count[14]), .Z(n32533)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_408.init = 16'heeee;
    LUT4 i1_2_lut_rep_296_3_lut (.A(count[15]), .B(count[14]), .C(n28430), 
         .Z(n32421)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_296_3_lut.init = 16'hfefe;
    LUT4 i2_2_lut_rep_345_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .D(count[13]), .Z(n32470)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_rep_345_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_362_3_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .Z(n32487)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_362_3_lut.init = 16'hfefe;
    LUT4 n28511_bdd_4_lut_25315 (.A(n28511), .B(count[9]), .C(n28382), 
         .D(n32447), .Z(n54)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A ((C+(D))+!B))) */ ;
    defparam n28511_bdd_4_lut_25315.init = 16'h002e;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1493_17 (.A0(count[15]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27350), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_17.INIT0 = 16'hd222;
    defparam add_1493_17.INIT1 = 16'h0000;
    defparam add_1493_17.INJECT1_0 = "NO";
    defparam add_1493_17.INJECT1_1 = "NO";
    CCU2D add_1493_15 (.A0(count[13]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32526), .C1(GND_net), .D1(GND_net), .CIN(n27349), 
          .COUT(n27350), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_15.INIT0 = 16'hd222;
    defparam add_1493_15.INIT1 = 16'hd222;
    defparam add_1493_15.INJECT1_0 = "NO";
    defparam add_1493_15.INJECT1_1 = "NO";
    CCU2D add_1493_13 (.A0(count[11]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32526), .C1(GND_net), .D1(GND_net), .CIN(n27348), 
          .COUT(n27349), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_13.INIT0 = 16'hd222;
    defparam add_1493_13.INIT1 = 16'hd222;
    defparam add_1493_13.INJECT1_0 = "NO";
    defparam add_1493_13.INJECT1_1 = "NO";
    CCU2D add_1493_11 (.A0(count[9]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32526), .C1(GND_net), .D1(GND_net), .CIN(n27347), 
          .COUT(n27348), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_11.INIT0 = 16'hd222;
    defparam add_1493_11.INIT1 = 16'hd222;
    defparam add_1493_11.INJECT1_0 = "NO";
    defparam add_1493_11.INJECT1_1 = "NO";
    CCU2D add_1493_9 (.A0(count[7]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32526), .C1(GND_net), .D1(GND_net), .CIN(n27346), 
          .COUT(n27347), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_9.INIT0 = 16'hd222;
    defparam add_1493_9.INIT1 = 16'hd222;
    defparam add_1493_9.INJECT1_0 = "NO";
    defparam add_1493_9.INJECT1_1 = "NO";
    CCU2D add_1493_7 (.A0(count[5]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32526), .C1(GND_net), .D1(GND_net), .CIN(n27345), 
          .COUT(n27346), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_7.INIT0 = 16'hd222;
    defparam add_1493_7.INIT1 = 16'hd222;
    defparam add_1493_7.INJECT1_0 = "NO";
    defparam add_1493_7.INJECT1_1 = "NO";
    CCU2D add_1493_5 (.A0(count[3]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32526), .C1(GND_net), .D1(GND_net), .CIN(n27344), 
          .COUT(n27345), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_5.INIT0 = 16'hd222;
    defparam add_1493_5.INIT1 = 16'hd222;
    defparam add_1493_5.INJECT1_0 = "NO";
    defparam add_1493_5.INJECT1_1 = "NO";
    CCU2D add_1493_3 (.A0(count[1]), .B0(n32526), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32526), .C1(GND_net), .D1(GND_net), .CIN(n27343), 
          .COUT(n27344), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_3.INIT0 = 16'hd222;
    defparam add_1493_3.INIT1 = 16'hd222;
    defparam add_1493_3.INJECT1_0 = "NO";
    defparam add_1493_3.INJECT1_1 = "NO";
    CCU2D add_1493_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30526), .B1(n1060), .C1(count[0]), .D1(n1048), .COUT(n27343), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_1.INIT0 = 16'hF000;
    defparam add_1493_1.INIT1 = 16'ha565;
    defparam add_1493_1.INJECT1_0 = "NO";
    defparam add_1493_1.INJECT1_1 = "NO";
    LUT4 i24675_4_lut (.A(n54), .B(n32524), .C(n30140), .D(n10), .Z(n30942)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i24675_4_lut.init = 16'h3323;
    CCU2D sub_61_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27638), 
          .S0(n943[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_9.INIT1 = 16'h0000;
    defparam sub_61_add_2_9.INJECT1_0 = "NO";
    defparam sub_61_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27637), 
          .COUT(n27638), .S0(n943[5]), .S1(n943[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_7.INJECT1_0 = "NO";
    defparam sub_61_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27636), 
          .COUT(n27637), .S0(n943[3]), .S1(n943[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_5.INJECT1_0 = "NO";
    defparam sub_61_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27635), 
          .COUT(n27636), .S0(n943[1]), .S1(n943[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_3.INJECT1_0 = "NO";
    defparam sub_61_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27635), 
          .S1(n943[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_1.INIT0 = 16'hF000;
    defparam sub_61_add_2_1.INIT1 = 16'h5555;
    defparam sub_61_add_2_1.INJECT1_0 = "NO";
    defparam sub_61_add_2_1.INJECT1_1 = "NO";
    LUT4 i7_4_lut (.A(n30737), .B(count[12]), .C(n12), .D(n11840), .Z(n14198)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i7_4_lut.init = 16'h0010;
    LUT4 i4_4_lut (.A(n28511), .B(n32375), .C(n28382), .D(count[9]), 
         .Z(n12)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i4_4_lut.init = 16'h0c88;
    LUT4 i14466_2_lut (.A(n943[1]), .B(n30140), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14466_2_lut.init = 16'h2222;
    LUT4 i14467_2_lut (.A(n943[2]), .B(n30140), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14467_2_lut.init = 16'h2222;
    LUT4 i14468_2_lut (.A(n943[3]), .B(n30140), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14468_2_lut.init = 16'h2222;
    LUT4 i14469_2_lut (.A(n943[4]), .B(n30140), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14469_2_lut.init = 16'h2222;
    LUT4 i14470_2_lut (.A(n943[5]), .B(n30140), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14470_2_lut.init = 16'h2222;
    LUT4 i14471_2_lut (.A(n943[6]), .B(n30140), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14471_2_lut.init = 16'h2222;
    LUT4 i14472_2_lut (.A(n943[7]), .B(n30140), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14472_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (n1039, debug_c_c, n28337, GND_net, n31041, 
            n32375, rc_ch7_c, \register[5] , n12031, n31025) /* synthesis syn_module_defined=1 */ ;
    output n1039;
    input debug_c_c;
    input n28337;
    input GND_net;
    output n31041;
    input n32375;
    input rc_ch7_c;
    output [7:0]\register[5] ;
    input n12031;
    output n31025;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n30521, n32445, n6, n32519, n32467, n32522, n4, n10, 
        n30134;
    wire [7:0]n934;
    wire [7:0]n43;
    
    wire n32468, n32418, n30541, n32521, n32518, n28495, n28336, 
        n32466, n30482, n12, n8, n32443, n54, n1045, n1033, 
        n11927, n28403, n6_adj_131, n28300, n4_adj_132, n28218, 
        n32481, n30540, n30522, n29821;
    wire [15:0]n116;
    
    wire n14177, n30187, n30706, n24, n27358, n27357, n27356, 
        n27355, n27354, n27353, n27352, n27351, n27642, n27641, 
        n27640, n27639;
    
    LUT4 i1_2_lut_rep_320_3_lut (.A(count[9]), .B(n30521), .C(count[8]), 
         .Z(n32445)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_320_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_342_4_lut (.A(count[3]), .B(n6), .C(n32519), .D(count[0]), 
         .Z(n32467)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_342_4_lut.init = 16'h8000;
    LUT4 i10_3_lut_4_lut_4_lut (.A(n32522), .B(n32467), .C(n4), .D(n32445), 
         .Z(n10)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i10_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut (.A(n30134), .B(n934[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_adj_237 (.A(n30134), .B(n934[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_237.init = 16'h4444;
    LUT4 i1_2_lut_adj_238 (.A(n30134), .B(n934[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_238.init = 16'h4444;
    LUT4 i1_2_lut_adj_239 (.A(n30134), .B(n934[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_239.init = 16'h4444;
    LUT4 i1_2_lut_adj_240 (.A(n30134), .B(n934[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_240.init = 16'h4444;
    LUT4 i1_2_lut_adj_241 (.A(n30134), .B(n934[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_241.init = 16'h4444;
    LUT4 i1_2_lut_adj_242 (.A(n30134), .B(n934[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_242.init = 16'h4444;
    LUT4 i1_3_lut_rep_293_4_lut (.A(count[8]), .B(n32468), .C(n4), .D(n32522), 
         .Z(n32418)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_3_lut_rep_293_4_lut.init = 16'hfeee;
    FD1P3IX valid_48 (.D(n30541), .SP(n28337), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1039));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i24774_4_lut (.A(n32521), .B(n32518), .C(n28495), .D(n28336), 
         .Z(n31041)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i24774_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n32466), .B(n30482), .C(n12), .D(n8), .Z(n28336)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    LUT4 i5_4_lut (.A(n32445), .B(n30521), .C(n32443), .D(n4), .Z(n12)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i5_4_lut.init = 16'h3222;
    LUT4 i1_2_lut_adj_243 (.A(n54), .B(n30134), .Z(n8)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_243.init = 16'h4444;
    LUT4 i1_4_lut_adj_244 (.A(count[4]), .B(count[5]), .C(count[3]), .D(n6), 
         .Z(n4)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_244.init = 16'hccc8;
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n32375), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1045));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1045), .SP(n32375), .CK(debug_c_c), .Q(n1033));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_245 (.A(n11927), .B(count[12]), .C(n32521), .D(count[13]), 
         .Z(n30521)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_4_lut_adj_245.init = 16'hfffe;
    LUT4 i1_2_lut_adj_246 (.A(count[11]), .B(count[10]), .Z(n11927)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_adj_246.init = 16'heeee;
    LUT4 i1_2_lut_adj_247 (.A(n1045), .B(n1033), .Z(n30482)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_247.init = 16'hbbbb;
    LUT4 i3_4_lut (.A(n28403), .B(n6_adj_131), .C(count[8]), .D(n32519), 
         .Z(n28300)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_4_lut.init = 16'hfefc;
    LUT4 i3_4_lut_adj_248 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n28403)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_248.init = 16'hfffe;
    LUT4 i2_2_lut_adj_249 (.A(count[6]), .B(count[7]), .Z(n6_adj_131)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut_adj_249.init = 16'heeee;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n11927), .D(n4_adj_132), 
         .Z(n28495)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_250 (.A(n32522), .B(count[9]), .C(n28218), .D(count[8]), 
         .Z(n4_adj_132)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_250.init = 16'heccc;
    LUT4 i2_4_lut_adj_251 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28218)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_251.init = 16'hfeee;
    LUT4 i1_4_lut_adj_252 (.A(n32468), .B(count[8]), .C(n32522), .D(n32481), 
         .Z(n30134)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_252.init = 16'hfbbb;
    LUT4 i5_2_lut_rep_393 (.A(n1033), .B(n1045), .Z(n32518)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_393.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1033), .B(n1045), .C(n28495), .D(n32521), 
         .Z(n30540)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_rep_394 (.A(count[4]), .B(count[5]), .Z(n32519)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_394.init = 16'h8888;
    LUT4 i3_3_lut_rep_356_4_lut (.A(count[4]), .B(count[5]), .C(n6), .D(count[3]), 
         .Z(n32481)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_3_lut_rep_356_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_396 (.A(count[15]), .B(count[14]), .Z(n32521)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_396.init = 16'heeee;
    LUT4 i1_2_lut_rep_397 (.A(count[6]), .B(count[7]), .Z(n32522)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_397.init = 16'h8888;
    LUT4 i1_2_lut_rep_318_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(n32481), 
         .D(count[0]), .Z(n32443)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_318_3_lut_4_lut.init = 16'h8000;
    LUT4 i24803_3_lut_3_lut_4_lut (.A(n32521), .B(n28495), .C(n32418), 
         .D(n30522), .Z(n30541)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i24803_3_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 n29821_bdd_4_lut_25330 (.A(n29821), .B(count[9]), .C(n28300), 
         .D(n30521), .Z(n54)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A ((C+(D))+!B))) */ ;
    defparam n29821_bdd_4_lut_25330.init = 16'h002e;
    LUT4 i14595_2_lut_rep_341 (.A(n28300), .B(count[9]), .Z(n32466)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14595_2_lut_rep_341.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(n28300), .B(count[9]), .C(n30521), .Z(n30522)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[0]), .B(n32481), .C(n32522), .D(count[8]), 
         .Z(n29821)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_343 (.A(count[9]), .B(n30521), .Z(n32468)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_343.init = 16'heeee;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    LUT4 i24758_4_lut (.A(n54), .B(n30482), .C(n30134), .D(n10), .Z(n31025)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i24758_4_lut.init = 16'h3323;
    LUT4 i3_4_lut_adj_253 (.A(n32521), .B(n30187), .C(n11927), .D(n32375), 
         .Z(n14177)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_253.init = 16'h0400;
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    LUT4 i4_4_lut (.A(n30706), .B(n24), .C(n1033), .D(n1045), .Z(n30187)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i4_4_lut.init = 16'h0040;
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    LUT4 i24349_2_lut (.A(count[13]), .B(count[12]), .Z(n30706)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24349_2_lut.init = 16'heeee;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    LUT4 i31_3_lut (.A(n29821), .B(n28300), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i31_3_lut.init = 16'h3a3a;
    CCU2D add_1489_17 (.A0(count[15]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27358), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_17.INIT0 = 16'hd222;
    defparam add_1489_17.INIT1 = 16'h0000;
    defparam add_1489_17.INJECT1_0 = "NO";
    defparam add_1489_17.INJECT1_1 = "NO";
    CCU2D add_1489_15 (.A0(count[13]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32518), .C1(GND_net), .D1(GND_net), .CIN(n27357), 
          .COUT(n27358), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_15.INIT0 = 16'hd222;
    defparam add_1489_15.INIT1 = 16'hd222;
    defparam add_1489_15.INJECT1_0 = "NO";
    defparam add_1489_15.INJECT1_1 = "NO";
    CCU2D add_1489_13 (.A0(count[11]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32518), .C1(GND_net), .D1(GND_net), .CIN(n27356), 
          .COUT(n27357), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_13.INIT0 = 16'hd222;
    defparam add_1489_13.INIT1 = 16'hd222;
    defparam add_1489_13.INJECT1_0 = "NO";
    defparam add_1489_13.INJECT1_1 = "NO";
    CCU2D add_1489_11 (.A0(count[9]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32518), .C1(GND_net), .D1(GND_net), .CIN(n27355), 
          .COUT(n27356), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_11.INIT0 = 16'hd222;
    defparam add_1489_11.INIT1 = 16'hd222;
    defparam add_1489_11.INJECT1_0 = "NO";
    defparam add_1489_11.INJECT1_1 = "NO";
    CCU2D add_1489_9 (.A0(count[7]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32518), .C1(GND_net), .D1(GND_net), .CIN(n27354), 
          .COUT(n27355), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_9.INIT0 = 16'hd222;
    defparam add_1489_9.INIT1 = 16'hd222;
    defparam add_1489_9.INJECT1_0 = "NO";
    defparam add_1489_9.INJECT1_1 = "NO";
    CCU2D add_1489_7 (.A0(count[5]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32518), .C1(GND_net), .D1(GND_net), .CIN(n27353), 
          .COUT(n27354), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_7.INIT0 = 16'hd222;
    defparam add_1489_7.INIT1 = 16'hd222;
    defparam add_1489_7.INJECT1_0 = "NO";
    defparam add_1489_7.INJECT1_1 = "NO";
    CCU2D add_1489_5 (.A0(count[3]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32518), .C1(GND_net), .D1(GND_net), .CIN(n27352), 
          .COUT(n27353), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_5.INIT0 = 16'hd222;
    defparam add_1489_5.INIT1 = 16'hd222;
    defparam add_1489_5.INJECT1_0 = "NO";
    defparam add_1489_5.INJECT1_1 = "NO";
    CCU2D add_1489_3 (.A0(count[1]), .B0(n32518), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32518), .C1(GND_net), .D1(GND_net), .CIN(n27351), 
          .COUT(n27352), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_3.INIT0 = 16'hd222;
    defparam add_1489_3.INIT1 = 16'hd222;
    defparam add_1489_3.INJECT1_0 = "NO";
    defparam add_1489_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_254 (.A(n30134), .B(n934[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_254.init = 16'h4444;
    CCU2D add_1489_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30540), .B1(n1045), .C1(count[0]), .D1(n1033), .COUT(n27351), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_1.INIT0 = 16'hF000;
    defparam add_1489_1.INIT1 = 16'ha565;
    defparam add_1489_1.INJECT1_0 = "NO";
    defparam add_1489_1.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27642), 
          .S0(n934[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_9.INIT1 = 16'h0000;
    defparam sub_60_add_2_9.INJECT1_0 = "NO";
    defparam sub_60_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27641), 
          .COUT(n27642), .S0(n934[5]), .S1(n934[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_7.INJECT1_0 = "NO";
    defparam sub_60_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27640), 
          .COUT(n27641), .S0(n934[3]), .S1(n934[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_5.INJECT1_0 = "NO";
    defparam sub_60_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27639), 
          .COUT(n27640), .S0(n934[1]), .S1(n934[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_3.INJECT1_0 = "NO";
    defparam sub_60_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27639), 
          .S1(n934[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_1.INIT0 = 16'hF000;
    defparam sub_60_add_2_1.INIT1 = 16'h5555;
    defparam sub_60_add_2_1.INJECT1_0 = "NO";
    defparam sub_60_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (\register[4] , debug_c_c, n11987, n32375, GND_net, 
            n34347, n31050, rc_ch4_c, n30958, n1024, n28331) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\register[4] ;
    input debug_c_c;
    input n11987;
    input n32375;
    input GND_net;
    input n34347;
    output n31050;
    input rc_ch4_c;
    output n30958;
    output n1024;
    input n28331;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n14143;
    wire [7:0]n43;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n30242, n32401, n18, n32384;
    wire [15:0]n116;
    
    wire n30185, n1018, n30598, n32427, n32426, n30441, n30490, 
        n28387, n1030, n30494, n32492, n32493, n30489, n32377, 
        n32410, n32402, n20339, n32458, n11813, n11779;
    wire [7:0]n925;
    
    wire n30459, n30741, n28407, n4, n30495, n32475, n6, n128_adj_129, 
        n5, n6_adj_130, n28404, n27366, n27365, n27364, n27363, 
        n27362, n27361, n27360, n27359, n27646, n27645, n27644, 
        n27643;
    
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_276 (.A(count[0]), .B(n30242), .Z(n32401)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_276.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[0]), .B(n30242), .C(count[9]), 
         .D(count[8]), .Z(n18)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf8f0;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_259_3_lut (.A(count[0]), .B(n30242), .C(count[8]), 
         .Z(n32384)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_259_3_lut.init = 16'h8080;
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(n32375), .B(n30185), .C(n1018), .D(n30598), .Z(n14143)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut.init = 16'h0080;
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    LUT4 i24797_3_lut_4_lut_4_lut (.A(n32427), .B(n30598), .C(n32426), 
         .D(n30441), .Z(n30490)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i24797_3_lut_4_lut_4_lut.init = 16'h1110;
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_226 (.A(n28387), .B(n1030), .C(n34347), .D(n18), 
         .Z(n30185)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_226.init = 16'h0200;
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(count[10]), .B(count[11]), .Z(n30494)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_367 (.A(n1030), .B(n1018), .Z(n32492)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_367.init = 16'hbbbb;
    LUT4 i24783_2_lut_3_lut (.A(n1030), .B(n1018), .C(n28387), .Z(n31050)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i24783_2_lut_3_lut.init = 16'h4040;
    LUT4 i5_2_lut_rep_368 (.A(n1018), .B(n1030), .Z(n32493)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_368.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n1018), .B(n1030), .C(n32427), .Z(n30489)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    FD1P3AX prev_in_46 (.D(n1030), .SP(n32375), .CK(debug_c_c), .Q(n1018));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n32375), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1030));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n32377), .B(n32410), .C(n32402), .D(n20339), .Z(n28387)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut.init = 16'heefe;
    LUT4 i21_3_lut_rep_252_4_lut (.A(count[8]), .B(n32401), .C(n32458), 
         .D(n30598), .Z(n32377)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21_3_lut_rep_252_4_lut.init = 16'h00f8;
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_227 (.A(count[15]), .B(count[14]), .Z(n11813)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_227.init = 16'heeee;
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_333 (.A(count[9]), .B(n11779), .Z(n32458)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_333.init = 16'heeee;
    LUT4 i1_3_lut_rep_285_4_lut (.A(count[9]), .B(n11779), .C(n30242), 
         .D(count[8]), .Z(n32410)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_3_lut_rep_285_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_301_3_lut (.A(count[9]), .B(n11779), .C(count[8]), 
         .Z(n32426)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_301_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_277_3_lut_4_lut (.A(count[9]), .B(n11779), .C(n30441), 
         .D(count[8]), .Z(n32402)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_277_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    LUT4 i14465_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14465_2_lut_4_lut.init = 16'h0200;
    LUT4 i24691_4_lut (.A(n30459), .B(n32493), .C(n32427), .D(n32492), 
         .Z(n30958)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i24691_4_lut.init = 16'h3031;
    LUT4 i3_4_lut_adj_228 (.A(n32426), .B(n30741), .C(n32401), .D(n30441), 
         .Z(n30459)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut_adj_228.init = 16'h3222;
    LUT4 i2_4_lut_adj_229 (.A(n30494), .B(count[9]), .C(n28407), .D(n4), 
         .Z(n30495)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_229.init = 16'hfeee;
    LUT4 i1_2_lut_3_lut_adj_230 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut_adj_230.init = 16'h8080;
    LUT4 i1_2_lut_rep_350_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), 
         .Z(n32475)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_350_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[2]), 
         .D(count[5]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_231 (.A(count[3]), .B(count[4]), .C(n128_adj_129), 
         .D(count[5]), .Z(n28407)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_231.init = 16'hffec;
    LUT4 i1_2_lut_adj_232 (.A(count[2]), .B(count[1]), .Z(n128_adj_129)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_232.init = 16'h8888;
    LUT4 i14257_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14257_2_lut_4_lut.init = 16'h0200;
    LUT4 i24244_4_lut (.A(n11779), .B(count[9]), .C(n5), .D(n6_adj_130), 
         .Z(n30598)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i24244_4_lut.init = 16'heeea;
    LUT4 i1_4_lut (.A(count[7]), .B(count[4]), .C(count[5]), .D(n28404), 
         .Z(n5)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_4_lut.init = 16'heaaa;
    LUT4 i2_2_lut (.A(count[8]), .B(count[6]), .Z(n6_adj_130)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_233 (.A(count[1]), .B(count[3]), .C(count[2]), .D(count[0]), 
         .Z(n28404)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_4_lut_adj_233.init = 16'hfffe;
    LUT4 i1_4_lut_adj_234 (.A(n128_adj_129), .B(n32475), .C(count[4]), 
         .D(count[3]), .Z(n30441)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_4_lut_adj_234.init = 16'hccc8;
    LUT4 i24383_3_lut_4_lut (.A(n32384), .B(n30598), .C(n32458), .D(n32410), 
         .Z(n30741)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i24383_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX valid_48 (.D(n30490), .SP(n28331), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1024));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_235 (.A(count[1]), .B(count[3]), .C(n6), .D(count[4]), 
         .Z(n30242)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_235.init = 16'h8000;
    CCU2D add_1485_17 (.A0(count[15]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27366), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_17.INIT0 = 16'hd222;
    defparam add_1485_17.INIT1 = 16'h0000;
    defparam add_1485_17.INJECT1_0 = "NO";
    defparam add_1485_17.INJECT1_1 = "NO";
    CCU2D add_1485_15 (.A0(count[13]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32493), .C1(GND_net), .D1(GND_net), .CIN(n27365), 
          .COUT(n27366), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_15.INIT0 = 16'hd222;
    defparam add_1485_15.INIT1 = 16'hd222;
    defparam add_1485_15.INJECT1_0 = "NO";
    defparam add_1485_15.INJECT1_1 = "NO";
    LUT4 i14601_2_lut_3_lut_4_lut (.A(count[8]), .B(n32458), .C(n30242), 
         .D(count[0]), .Z(n20339)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i14601_2_lut_3_lut_4_lut.init = 16'hfeee;
    CCU2D add_1485_13 (.A0(count[11]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32493), .C1(GND_net), .D1(GND_net), .CIN(n27364), 
          .COUT(n27365), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_13.INIT0 = 16'hd222;
    defparam add_1485_13.INIT1 = 16'hd222;
    defparam add_1485_13.INJECT1_0 = "NO";
    defparam add_1485_13.INJECT1_1 = "NO";
    CCU2D add_1485_11 (.A0(count[9]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32493), .C1(GND_net), .D1(GND_net), .CIN(n27363), 
          .COUT(n27364), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_11.INIT0 = 16'hd222;
    defparam add_1485_11.INIT1 = 16'hd222;
    defparam add_1485_11.INJECT1_0 = "NO";
    defparam add_1485_11.INJECT1_1 = "NO";
    CCU2D add_1485_9 (.A0(count[7]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32493), .C1(GND_net), .D1(GND_net), .CIN(n27362), 
          .COUT(n27363), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_9.INIT0 = 16'hd222;
    defparam add_1485_9.INIT1 = 16'hd222;
    defparam add_1485_9.INJECT1_0 = "NO";
    defparam add_1485_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_302 (.A(n11813), .B(count[13]), .C(count[12]), .D(n30495), 
         .Z(n32427)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_302.init = 16'heaaa;
    CCU2D add_1485_7 (.A0(count[5]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32493), .C1(GND_net), .D1(GND_net), .CIN(n27361), 
          .COUT(n27362), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_7.INIT0 = 16'hd222;
    defparam add_1485_7.INIT1 = 16'hd222;
    defparam add_1485_7.INJECT1_0 = "NO";
    defparam add_1485_7.INJECT1_1 = "NO";
    CCU2D add_1485_5 (.A0(count[3]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32493), .C1(GND_net), .D1(GND_net), .CIN(n27360), 
          .COUT(n27361), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_5.INIT0 = 16'hd222;
    defparam add_1485_5.INIT1 = 16'hd222;
    defparam add_1485_5.INJECT1_0 = "NO";
    defparam add_1485_5.INJECT1_1 = "NO";
    CCU2D add_1485_3 (.A0(count[1]), .B0(n32493), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32493), .C1(GND_net), .D1(GND_net), .CIN(n27359), 
          .COUT(n27360), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_3.INIT0 = 16'hd222;
    defparam add_1485_3.INIT1 = 16'hd222;
    defparam add_1485_3.INJECT1_0 = "NO";
    defparam add_1485_3.INJECT1_1 = "NO";
    CCU2D add_1485_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30489), .B1(n1030), .C1(count[0]), .D1(n1018), .COUT(n27359), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_1.INIT0 = 16'hF000;
    defparam add_1485_1.INIT1 = 16'ha565;
    defparam add_1485_1.INJECT1_0 = "NO";
    defparam add_1485_1.INJECT1_1 = "NO";
    LUT4 i14459_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14459_2_lut_4_lut.init = 16'h0200;
    LUT4 i14460_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14460_2_lut_4_lut.init = 16'h0200;
    CCU2D sub_59_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27646), 
          .S0(n925[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_9.INIT1 = 16'h0000;
    defparam sub_59_add_2_9.INJECT1_0 = "NO";
    defparam sub_59_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27645), 
          .COUT(n27646), .S0(n925[5]), .S1(n925[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_7.INJECT1_0 = "NO";
    defparam sub_59_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27644), 
          .COUT(n27645), .S0(n925[3]), .S1(n925[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_5.INJECT1_0 = "NO";
    defparam sub_59_add_2_5.INJECT1_1 = "NO";
    LUT4 i14462_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14462_2_lut_4_lut.init = 16'h0200;
    CCU2D sub_59_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27643), 
          .COUT(n27644), .S0(n925[1]), .S1(n925[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_3.INJECT1_0 = "NO";
    defparam sub_59_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27643), 
          .S1(n925[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_1.INIT0 = 16'hF000;
    defparam sub_59_add_2_1.INIT1 = 16'h5555;
    defparam sub_59_add_2_1.INJECT1_0 = "NO";
    defparam sub_59_add_2_1.INJECT1_1 = "NO";
    LUT4 i14463_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14463_2_lut_4_lut.init = 16'h0200;
    LUT4 i14461_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14461_2_lut_4_lut.init = 16'h0200;
    LUT4 i3_4_lut_adj_236 (.A(count[12]), .B(count[13]), .C(n11813), .D(n30494), 
         .Z(n11779)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_236.init = 16'hfffe;
    LUT4 i14464_2_lut_4_lut (.A(count[8]), .B(n30242), .C(n32458), .D(n925[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14464_2_lut_4_lut.init = 16'h0200;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (debug_c_c, n32375, GND_net, \register[3] , n12138, 
            n1009, n28345, n30999, rc_ch3_c, n31033) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n32375;
    input GND_net;
    output [7:0]\register[3] ;
    input n12138;
    output n1009;
    input n28345;
    output n30999;
    input rc_ch3_c;
    output n31033;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    wire [15:0]n116;
    
    wire n152, n103, n154, n32531, n32532, n6, n14451;
    wire [7:0]n43;
    
    wire n32517, n32516, n32464, n32465;
    wire [7:0]n916;
    
    wire n54, n7, n30544, n30515, n32444, n10, n32520, n11, 
        n30765, n26, n1003, n1015, n30466, n4, n28208, n32515, 
        n11819, n32514, n28497, n28343, n5, n20343, n6_adj_126, 
        n30581, n4_adj_127, n32479, n4_adj_128, n30543, n32417, 
        n32480, n27370, n27371, n27369, n27368, n27367, n27374, 
        n27373, n27650, n27372, n27649, n27648, n27647;
    
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    PFUMX i13432 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    LUT4 i23_4_lut (.A(n32531), .B(count[2]), .C(n32532), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    LUT4 i3_3_lut_rep_339_4_lut (.A(count[3]), .B(n32532), .C(n32517), 
         .D(n32516), .Z(n32464)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_3_lut_rep_339_4_lut.init = 16'h8000;
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i14455_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14455_2_lut_4_lut.init = 16'h0400;
    LUT4 i14454_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14454_2_lut_4_lut.init = 16'h0400;
    LUT4 i14453_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14453_2_lut_4_lut.init = 16'h0400;
    LUT4 i14452_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14452_2_lut_4_lut.init = 16'h0400;
    LUT4 i14451_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14451_2_lut_4_lut.init = 16'h0400;
    LUT4 i14450_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14450_2_lut_4_lut.init = 16'h0400;
    LUT4 i14449_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14449_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n54), 
         .Z(n7)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h00fb;
    LUT4 i14252_2_lut_4_lut (.A(n32465), .B(count[8]), .C(n32464), .D(n916[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14252_2_lut_4_lut.init = 16'h0400;
    FD1P3IX valid_48 (.D(n30544), .SP(n28345), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1009));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i24732_4_lut (.A(n54), .B(n30515), .C(n32444), .D(n10), .Z(n30999)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i24732_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n32375), .B(n32520), .C(n11), .D(n30765), .Z(n14451)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i4_3_lut (.A(n26), .B(n1003), .C(n1015), .Z(n11)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i4_3_lut.init = 16'h0808;
    LUT4 i33_4_lut (.A(count[8]), .B(n154), .C(count[9]), .D(n30466), 
         .Z(n26)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i33_4_lut.init = 16'h3a30;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n32375), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1015));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1015), .SP(n32375), .CK(debug_c_c), .Q(n1003));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_220 (.A(n32517), .B(count[5]), .C(count[3]), .D(n4), 
         .Z(n28208)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_220.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n32520), .D(n32515), 
         .Z(n11819)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i24766_4_lut (.A(n32520), .B(n32514), .C(n28497), .D(n28343), 
         .Z(n31033)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i24766_4_lut.init = 16'h3233;
    LUT4 i21_4_lut (.A(n5), .B(n20343), .C(n32465), .D(n6_adj_126), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_4_lut (.A(n20343), .B(n30515), .C(n7), .D(n30581), .Z(n28343)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    LUT4 i1_2_lut (.A(n1015), .B(n1003), .Z(n30515)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i14605_3_lut (.A(count[9]), .B(n11819), .C(n154), .Z(n20343)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i14605_3_lut.init = 16'hecec;
    LUT4 i2_4_lut_adj_221 (.A(count[13]), .B(count[12]), .C(n32515), .D(n4_adj_127), 
         .Z(n28497)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_221.init = 16'h8880;
    LUT4 i1_4_lut_adj_222 (.A(count[9]), .B(count[4]), .C(n32479), .D(n4_adj_128), 
         .Z(n4_adj_127)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_222.init = 16'hfaea;
    LUT4 i5_2_lut_rep_389 (.A(n1003), .B(n1015), .Z(n32514)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_389.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1003), .B(n1015), .C(n28497), .D(n32520), 
         .Z(n30543)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_rep_390 (.A(count[10]), .B(count[11]), .Z(n32515)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_390.init = 16'heeee;
    LUT4 i24407_3_lut_4_lut (.A(count[10]), .B(count[11]), .C(count[13]), 
         .D(count[12]), .Z(n30765)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24407_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_391 (.A(count[2]), .B(count[1]), .Z(n32516)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_391.init = 16'h8888;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(n32517), 
         .D(count[8]), .Z(n6_adj_126)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4_adj_128)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_392 (.A(count[6]), .B(count[7]), .Z(n32517)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_392.init = 16'h8888;
    LUT4 i1_2_lut_rep_354_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n32479)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_354_3_lut.init = 16'h8080;
    LUT4 i24795_3_lut_3_lut_4_lut (.A(n32520), .B(n28497), .C(n32417), 
         .D(n20343), .Z(n30544)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i24795_3_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_395 (.A(count[15]), .B(count[14]), .Z(n32520)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_395.init = 16'heeee;
    LUT4 i2_3_lut_rep_406 (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n32531)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_406.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_223 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .D(n32532), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_223.init = 16'hfffe;
    LUT4 i1_2_lut_rep_407 (.A(count[4]), .B(count[5]), .Z(n32532)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_407.init = 16'h8888;
    LUT4 i1_2_lut_rep_355_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n32480)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_355_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_224 (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n5)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut_4_lut_adj_224.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_225 (.A(n32516), .B(n32517), .C(n32480), .D(count[0]), 
         .Z(n30466)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_225.init = 16'h8000;
    LUT4 i1_2_lut_rep_340 (.A(count[9]), .B(n11819), .Z(n32465)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_340.init = 16'heeee;
    LUT4 i1_2_lut_rep_292_3_lut_4_lut (.A(count[9]), .B(n11819), .C(n28208), 
         .D(count[8]), .Z(n32417)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_292_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_rep_319_4_lut (.A(count[9]), .B(n11819), .C(n32464), 
         .D(count[8]), .Z(n32444)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_3_lut_rep_319_4_lut.init = 16'hfeff;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n32465), .C(n30466), 
         .D(n28208), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i24229_3_lut_4_lut (.A(count[8]), .B(n32465), .C(n28208), .D(n30466), 
         .Z(n30581)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i24229_3_lut_4_lut.init = 16'hfeee;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1481_9 (.A0(count[7]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32514), .C1(GND_net), .D1(GND_net), .CIN(n27370), 
          .COUT(n27371), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_9.INIT0 = 16'hd222;
    defparam add_1481_9.INIT1 = 16'hd222;
    defparam add_1481_9.INJECT1_0 = "NO";
    defparam add_1481_9.INJECT1_1 = "NO";
    CCU2D add_1481_7 (.A0(count[5]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32514), .C1(GND_net), .D1(GND_net), .CIN(n27369), 
          .COUT(n27370), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_7.INIT0 = 16'hd222;
    defparam add_1481_7.INIT1 = 16'hd222;
    defparam add_1481_7.INJECT1_0 = "NO";
    defparam add_1481_7.INJECT1_1 = "NO";
    CCU2D add_1481_5 (.A0(count[3]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32514), .C1(GND_net), .D1(GND_net), .CIN(n27368), 
          .COUT(n27369), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_5.INIT0 = 16'hd222;
    defparam add_1481_5.INIT1 = 16'hd222;
    defparam add_1481_5.INJECT1_0 = "NO";
    defparam add_1481_5.INJECT1_1 = "NO";
    CCU2D add_1481_3 (.A0(count[1]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32514), .C1(GND_net), .D1(GND_net), .CIN(n27367), 
          .COUT(n27368), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_3.INIT0 = 16'hd222;
    defparam add_1481_3.INIT1 = 16'hd222;
    defparam add_1481_3.INJECT1_0 = "NO";
    defparam add_1481_3.INJECT1_1 = "NO";
    CCU2D add_1481_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30543), .B1(n1015), .C1(count[0]), .D1(n1003), .COUT(n27367), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_1.INIT0 = 16'hF000;
    defparam add_1481_1.INIT1 = 16'ha565;
    defparam add_1481_1.INJECT1_0 = "NO";
    defparam add_1481_1.INJECT1_1 = "NO";
    CCU2D add_1481_17 (.A0(count[15]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27374), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_17.INIT0 = 16'hd222;
    defparam add_1481_17.INIT1 = 16'h0000;
    defparam add_1481_17.INJECT1_0 = "NO";
    defparam add_1481_17.INJECT1_1 = "NO";
    CCU2D add_1481_15 (.A0(count[13]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32514), .C1(GND_net), .D1(GND_net), .CIN(n27373), 
          .COUT(n27374), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_15.INIT0 = 16'hd222;
    defparam add_1481_15.INIT1 = 16'hd222;
    defparam add_1481_15.INJECT1_0 = "NO";
    defparam add_1481_15.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27650), 
          .S0(n916[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_9.INIT1 = 16'h0000;
    defparam sub_58_add_2_9.INJECT1_0 = "NO";
    defparam sub_58_add_2_9.INJECT1_1 = "NO";
    CCU2D add_1481_13 (.A0(count[11]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32514), .C1(GND_net), .D1(GND_net), .CIN(n27372), 
          .COUT(n27373), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_13.INIT0 = 16'hd222;
    defparam add_1481_13.INIT1 = 16'hd222;
    defparam add_1481_13.INJECT1_0 = "NO";
    defparam add_1481_13.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27649), 
          .COUT(n27650), .S0(n916[5]), .S1(n916[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_7.INJECT1_0 = "NO";
    defparam sub_58_add_2_7.INJECT1_1 = "NO";
    CCU2D add_1481_11 (.A0(count[9]), .B0(n32514), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32514), .C1(GND_net), .D1(GND_net), .CIN(n27371), 
          .COUT(n27372), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_11.INIT0 = 16'hd222;
    defparam add_1481_11.INIT1 = 16'hd222;
    defparam add_1481_11.INJECT1_0 = "NO";
    defparam add_1481_11.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27648), 
          .COUT(n27649), .S0(n916[3]), .S1(n916[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_5.INJECT1_0 = "NO";
    defparam sub_58_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27647), 
          .COUT(n27648), .S0(n916[1]), .S1(n916[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_3.INJECT1_0 = "NO";
    defparam sub_58_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27647), 
          .S1(n916[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_1.INIT0 = 16'hF000;
    defparam sub_58_add_2_1.INIT1 = 16'h5555;
    defparam sub_58_add_2_1.INJECT1_0 = "NO";
    defparam sub_58_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (debug_c_c, n32375, GND_net, \register[2] , n32369, 
            n14446, n994, n1000, n988, rc_ch2_c, n54, n4) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n32375;
    input GND_net;
    output [7:0]\register[2] ;
    input n32369;
    input n14446;
    output n994;
    output n1000;
    output n988;
    input rc_ch2_c;
    output n54;
    output n4;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n32541, n28281, n4_c;
    wire [15:0]n116;
    wire [7:0]n43;
    
    wire n30289, n11825, n32549, n30343, n29754, n32548, n28223, 
        n30465, n30464, n28088, n32496, n4_adj_123, n5, n30675, 
        n20403, n8, n32366, n30485, n32540, n63, n21791, n30546, 
        n30767, n25, n11, n6, n4_adj_124, n32456, n32455, n32476, 
        n27382, n27381, n27380, n27379, n27378, n27377, n27376, 
        n27375, n27654;
    wire [7:0]n907;
    
    wire n27653, n27652, n27651, n29825, n28411;
    
    LUT4 i1_3_lut_4_lut (.A(count[8]), .B(n32541), .C(count[9]), .D(n28281), 
         .Z(n4_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i1_4_lut_then_4_lut (.A(n30289), .B(n11825), .C(count[9]), .D(n32541), 
         .Z(n32549)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+(C)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0103;
    LUT4 i1_4_lut_else_4_lut (.A(n30343), .B(n29754), .C(n11825), .D(count[9]), 
         .Z(n32548)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0002;
    FD1P3AX valid_48 (.D(n30465), .SP(n28223), .CK(debug_c_c), .Q(n994));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i24787_4_lut (.A(n1000), .B(n30464), .C(n988), .D(n32375), 
         .Z(n28223)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(D)))) */ ;
    defparam i24787_4_lut.init = 16'h3100;
    LUT4 i1_4_lut (.A(n28088), .B(n32496), .C(n988), .D(n4_adj_123), 
         .Z(n30464)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h1101;
    LUT4 i1_4_lut_adj_201 (.A(n1000), .B(n5), .C(n30675), .D(n20403), 
         .Z(n4_adj_123)) /* synthesis lut_function=(A+!(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_201.init = 16'haaea;
    LUT4 i2_4_lut (.A(n32496), .B(count[12]), .C(n8), .D(count[11]), 
         .Z(n30465)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut.init = 16'h0010;
    LUT4 i3_3_lut (.A(n32366), .B(count[10]), .C(count[13]), .Z(n8)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i3_3_lut.init = 16'h0202;
    LUT4 i2_4_lut_adj_202 (.A(count[12]), .B(n30485), .C(count[13]), .D(n4_c), 
         .Z(n28088)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_202.init = 16'ha080;
    LUT4 i2_4_lut_adj_203 (.A(count[3]), .B(count[5]), .C(n32540), .D(count[4]), 
         .Z(n28281)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_203.init = 16'hffec;
    LUT4 i1_2_lut (.A(n1000), .B(n988), .Z(n63)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_adj_204 (.A(n1000), .B(n988), .Z(n21791)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_204.init = 16'h2222;
    LUT4 i1_2_lut_rep_371 (.A(count[14]), .B(count[15]), .Z(n32496)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_371.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[14]), .B(count[15]), .C(n21791), .D(n28088), 
         .Z(n30546)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 count_8__bdd_4_lut (.A(count[8]), .B(n30343), .C(n30767), .D(count[9]), 
         .Z(n32366)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam count_8__bdd_4_lut.init = 16'hf0ee;
    LUT4 i24840_4_lut (.A(count[8]), .B(count[7]), .C(n25), .D(count[6]), 
         .Z(n30767)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24840_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_205 (.A(count[0]), .B(n11), .C(n6), .D(count[1]), 
         .Z(n25)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_205.init = 16'hccc8;
    LUT4 i2_2_lut (.A(count[3]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_206 (.A(n32541), .B(count[5]), .C(count[4]), .D(n4_adj_124), 
         .Z(n30343)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_206.init = 16'h8880;
    LUT4 i1_2_lut_adj_207 (.A(count[5]), .B(count[4]), .Z(n11)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_207.init = 16'h8888;
    LUT4 i1_2_lut_rep_331 (.A(count[9]), .B(n11825), .Z(n32456)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_331.init = 16'heeee;
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n32375), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1000));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1000), .SP(n32375), .CK(debug_c_c), .Q(n988));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_415 (.A(count[2]), .B(count[1]), .Z(n32540)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_415.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[3]), .Z(n4_adj_124)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_416 (.A(count[6]), .B(count[7]), .Z(n32541)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_416.init = 16'h8888;
    LUT4 i1_2_lut_rep_330_3_lut (.A(count[6]), .B(count[7]), .C(n30289), 
         .Z(n32455)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_330_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[0]), 
         .D(n30289), .Z(n29754)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_351_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n32476)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_351_3_lut.init = 16'h8080;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n32369), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1477_17 (.A0(count[15]), .B0(n63), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27382), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_17.INIT0 = 16'h7888;
    defparam add_1477_17.INIT1 = 16'h0000;
    defparam add_1477_17.INJECT1_0 = "NO";
    defparam add_1477_17.INJECT1_1 = "NO";
    CCU2D add_1477_15 (.A0(n63), .B0(count[13]), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n63), .C1(GND_net), .D1(GND_net), .CIN(n27381), 
          .COUT(n27382), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_15.INIT0 = 16'h7888;
    defparam add_1477_15.INIT1 = 16'h7888;
    defparam add_1477_15.INJECT1_0 = "NO";
    defparam add_1477_15.INJECT1_1 = "NO";
    CCU2D add_1477_13 (.A0(count[11]), .B0(n21791), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n63), .C1(GND_net), .D1(GND_net), .CIN(n27380), 
          .COUT(n27381), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_13.INIT0 = 16'hd222;
    defparam add_1477_13.INIT1 = 16'h7888;
    defparam add_1477_13.INJECT1_0 = "NO";
    defparam add_1477_13.INJECT1_1 = "NO";
    CCU2D add_1477_11 (.A0(count[9]), .B0(n21791), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n21791), .C1(GND_net), .D1(GND_net), .CIN(n27379), 
          .COUT(n27380), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_11.INIT0 = 16'hd222;
    defparam add_1477_11.INIT1 = 16'hd222;
    defparam add_1477_11.INJECT1_0 = "NO";
    defparam add_1477_11.INJECT1_1 = "NO";
    CCU2D add_1477_9 (.A0(count[7]), .B0(n21791), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n21791), .C1(GND_net), .D1(GND_net), .CIN(n27378), 
          .COUT(n27379), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_9.INIT0 = 16'hd222;
    defparam add_1477_9.INIT1 = 16'hd222;
    defparam add_1477_9.INJECT1_0 = "NO";
    defparam add_1477_9.INJECT1_1 = "NO";
    CCU2D add_1477_7 (.A0(count[5]), .B0(n21791), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n21791), .C1(GND_net), .D1(GND_net), .CIN(n27377), 
          .COUT(n27378), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_7.INIT0 = 16'hd222;
    defparam add_1477_7.INIT1 = 16'hd222;
    defparam add_1477_7.INJECT1_0 = "NO";
    defparam add_1477_7.INJECT1_1 = "NO";
    CCU2D add_1477_5 (.A0(count[3]), .B0(n21791), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n21791), .C1(GND_net), .D1(GND_net), .CIN(n27376), 
          .COUT(n27377), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_5.INIT0 = 16'hd222;
    defparam add_1477_5.INIT1 = 16'hd222;
    defparam add_1477_5.INJECT1_0 = "NO";
    defparam add_1477_5.INJECT1_1 = "NO";
    CCU2D add_1477_3 (.A0(count[1]), .B0(n21791), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n21791), .C1(GND_net), .D1(GND_net), .CIN(n27375), 
          .COUT(n27376), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_3.INIT0 = 16'hd222;
    defparam add_1477_3.INIT1 = 16'hd222;
    defparam add_1477_3.INJECT1_0 = "NO";
    defparam add_1477_3.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27654), 
          .S0(n907[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_9.INIT1 = 16'h0000;
    defparam sub_57_add_2_9.INJECT1_0 = "NO";
    defparam sub_57_add_2_9.INJECT1_1 = "NO";
    CCU2D add_1477_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30546), .B1(n1000), .C1(count[0]), .D1(n988), .COUT(n27375), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_1.INIT0 = 16'hF000;
    defparam add_1477_1.INIT1 = 16'ha565;
    defparam add_1477_1.INJECT1_0 = "NO";
    defparam add_1477_1.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27653), 
          .COUT(n27654), .S0(n907[5]), .S1(n907[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_7.INJECT1_0 = "NO";
    defparam sub_57_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27652), 
          .COUT(n27653), .S0(n907[3]), .S1(n907[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_5.INJECT1_0 = "NO";
    defparam sub_57_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27651), 
          .COUT(n27652), .S0(n907[1]), .S1(n907[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_3.INJECT1_0 = "NO";
    defparam sub_57_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27651), 
          .S1(n907[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_1.INIT0 = 16'hF000;
    defparam sub_57_add_2_1.INIT1 = 16'h5555;
    defparam sub_57_add_2_1.INJECT1_0 = "NO";
    defparam sub_57_add_2_1.INJECT1_1 = "NO";
    LUT4 i24320_3_lut_4_lut (.A(count[8]), .B(n32456), .C(n30343), .D(n29754), 
         .Z(n30675)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i24320_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_4_lut (.A(n32455), .B(count[8]), .C(n32456), .D(n907[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_208 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n54), .Z(n5)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_208.init = 16'h00fb;
    LUT4 i21_4_lut (.A(n29825), .B(n20403), .C(n32456), .D(n32476), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_2_lut_adj_209 (.A(count[0]), .B(n30289), .Z(n29825)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_209.init = 16'h8888;
    LUT4 i3_4_lut (.A(count[3]), .B(n11), .C(count[1]), .D(count[2]), 
         .Z(n30289)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_210 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n907[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_210.init = 16'h0400;
    LUT4 i14665_3_lut (.A(n28411), .B(n11825), .C(count[9]), .Z(n20403)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i14665_3_lut.init = 16'hecec;
    LUT4 i3_4_lut_adj_211 (.A(n25), .B(count[6]), .C(count[8]), .D(count[7]), 
         .Z(n28411)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_211.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_212 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n907[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_212.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_213 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n907[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_213.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_214 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n907[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_214.init = 16'h0400;
    LUT4 i3_4_lut_adj_215 (.A(count[13]), .B(n30485), .C(count[12]), .D(n32496), 
         .Z(n11825)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_215.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_216 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n907[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_216.init = 16'h0400;
    LUT4 i1_2_lut_adj_217 (.A(count[10]), .B(count[11]), .Z(n30485)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_217.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_218 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n907[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_218.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_219 (.A(n32455), .B(count[8]), .C(n32456), 
         .D(n907[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_219.init = 16'h0400;
    PFUMX i25283 (.BLUT(n32548), .ALUT(n32549), .C0(count[8]), .Z(n4));
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (debug_c_c, n32375, GND_net, \register[1] , n32374, 
            n31079, n979, n28339, rc_ch1_c, n30940) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n32375;
    input GND_net;
    output [7:0]\register[1] ;
    input n32374;
    output n31079;
    output n979;
    input n28339;
    input rc_ch1_c;
    output n30940;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    wire [15:0]n116;
    
    wire n14448;
    wire [7:0]n43;
    
    wire n30353, n32434, n30668, n32433, n30504, n54, n973, n985, 
        n32497, n30505, n4, n30352, n11792, n32457, n27390, n30548, 
        n23, n10;
    wire [7:0]n898;
    
    wire n27389, n30347, n95, n27388, n27387, n27386, n27385, 
        n11845, n30527, n27384, n27383, n27658, n27657, n27656, 
        n6, n27655, n49_adj_122, n30781, n30745, n30170, n30761, 
        n28414, n30529;
    
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i24680_3_lut_3_lut_4_lut (.A(n30353), .B(n32434), .C(n30668), 
         .D(n32433), .Z(n30504)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i24680_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i8682_2_lut_3_lut (.A(n32375), .B(n31079), .C(n54), .Z(n14448)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i8682_2_lut_3_lut.init = 16'h8080;
    LUT4 i5_2_lut_rep_372 (.A(n973), .B(n985), .Z(n32497)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_372.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n973), .B(n985), .C(n32433), .Z(n30505)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_3_lut_adj_192 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut_adj_192.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_193 (.A(count[6]), .B(count[7]), .C(count[5]), 
         .Z(n30352)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut_adj_193.init = 16'h8080;
    LUT4 i1_2_lut_rep_332 (.A(count[9]), .B(n11792), .Z(n32457)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_332.init = 16'heeee;
    LUT4 i1_2_lut_rep_309_3_lut (.A(count[9]), .B(n11792), .C(count[8]), 
         .Z(n32434)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_309_3_lut.init = 16'hfefe;
    FD1P3AX valid_48 (.D(n30504), .SP(n28339), .CK(debug_c_c), .Q(n979));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n985), .SP(n32375), .CK(debug_c_c), .Q(n973));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n32375), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n985));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32375), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32375), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n32374), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1473_17 (.A0(count[15]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27390), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_17.INIT0 = 16'hd222;
    defparam add_1473_17.INIT1 = 16'h0000;
    defparam add_1473_17.INJECT1_0 = "NO";
    defparam add_1473_17.INJECT1_1 = "NO";
    LUT4 i24812_4_lut (.A(n54), .B(n30548), .C(n23), .D(n10), .Z(n31079)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i24812_4_lut.init = 16'h3332;
    LUT4 i14244_2_lut (.A(n898[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14244_2_lut.init = 16'h8888;
    CCU2D add_1473_15 (.A0(count[13]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32497), .C1(GND_net), .D1(GND_net), .CIN(n27389), 
          .COUT(n27390), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_15.INIT0 = 16'hd222;
    defparam add_1473_15.INIT1 = 16'hd222;
    defparam add_1473_15.INJECT1_0 = "NO";
    defparam add_1473_15.INJECT1_1 = "NO";
    LUT4 i21_4_lut (.A(count[8]), .B(n30668), .C(n32457), .D(n30347), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_2_lut (.A(n985), .B(n973), .Z(n30548)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut (.A(count[8]), .B(n32457), .C(count[1]), .D(n95), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0222;
    CCU2D add_1473_13 (.A0(count[11]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32497), .C1(GND_net), .D1(GND_net), .CIN(n27388), 
          .COUT(n27389), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_13.INIT0 = 16'hd222;
    defparam add_1473_13.INIT1 = 16'hd222;
    defparam add_1473_13.INJECT1_0 = "NO";
    defparam add_1473_13.INJECT1_1 = "NO";
    CCU2D add_1473_11 (.A0(count[9]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32497), .C1(GND_net), .D1(GND_net), .CIN(n27387), 
          .COUT(n27388), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_11.INIT0 = 16'hd222;
    defparam add_1473_11.INIT1 = 16'hd222;
    defparam add_1473_11.INJECT1_0 = "NO";
    defparam add_1473_11.INJECT1_1 = "NO";
    CCU2D add_1473_9 (.A0(count[7]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32497), .C1(GND_net), .D1(GND_net), .CIN(n27386), 
          .COUT(n27387), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_9.INIT0 = 16'hd222;
    defparam add_1473_9.INIT1 = 16'hd222;
    defparam add_1473_9.INJECT1_0 = "NO";
    defparam add_1473_9.INJECT1_1 = "NO";
    LUT4 i3_4_lut (.A(count[3]), .B(count[4]), .C(count[2]), .D(n30352), 
         .Z(n95)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut.init = 16'h8000;
    CCU2D add_1473_7 (.A0(count[5]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32497), .C1(GND_net), .D1(GND_net), .CIN(n27385), 
          .COUT(n27386), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_7.INIT0 = 16'hd222;
    defparam add_1473_7.INIT1 = 16'hd222;
    defparam add_1473_7.INJECT1_0 = "NO";
    defparam add_1473_7.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_194 (.A(count[12]), .B(count[13]), .C(n11845), .D(n30527), 
         .Z(n11792)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_194.init = 16'hfffe;
    LUT4 i1_2_lut_adj_195 (.A(count[15]), .B(count[14]), .Z(n11845)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_195.init = 16'heeee;
    CCU2D add_1473_5 (.A0(count[3]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32497), .C1(GND_net), .D1(GND_net), .CIN(n27384), 
          .COUT(n27385), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_5.INIT0 = 16'hd222;
    defparam add_1473_5.INIT1 = 16'hd222;
    defparam add_1473_5.INJECT1_0 = "NO";
    defparam add_1473_5.INJECT1_1 = "NO";
    CCU2D add_1473_3 (.A0(count[1]), .B0(n32497), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32497), .C1(GND_net), .D1(GND_net), .CIN(n27383), 
          .COUT(n27384), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_3.INIT0 = 16'hd222;
    defparam add_1473_3.INIT1 = 16'hd222;
    defparam add_1473_3.INJECT1_0 = "NO";
    defparam add_1473_3.INJECT1_1 = "NO";
    CCU2D add_1473_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30505), .B1(n985), .C1(count[0]), .D1(n973), .COUT(n27383), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_1.INIT0 = 16'hF000;
    defparam add_1473_1.INIT1 = 16'ha565;
    defparam add_1473_1.INJECT1_0 = "NO";
    defparam add_1473_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_196 (.A(count[11]), .B(count[10]), .Z(n30527)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_196.init = 16'heeee;
    LUT4 i2_3_lut (.A(n95), .B(count[1]), .C(count[0]), .Z(n30347)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_3_lut.init = 16'h8080;
    CCU2D sub_56_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27658), 
          .S0(n898[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_9.INIT1 = 16'h0000;
    defparam sub_56_add_2_9.INJECT1_0 = "NO";
    defparam sub_56_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27657), 
          .COUT(n27658), .S0(n898[5]), .S1(n898[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_7.INJECT1_0 = "NO";
    defparam sub_56_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27656), 
          .COUT(n27657), .S0(n898[3]), .S1(n898[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_5.INJECT1_0 = "NO";
    defparam sub_56_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_197 (.A(count[4]), .B(n30352), .C(count[3]), .D(n6), 
         .Z(n30353)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_4_lut_adj_197.init = 16'hccc8;
    CCU2D sub_56_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27655), 
          .COUT(n27656), .S0(n898[1]), .S1(n898[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_3.INJECT1_0 = "NO";
    defparam sub_56_add_2_3.INJECT1_1 = "NO";
    LUT4 i2786_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2786_2_lut.init = 16'h8888;
    CCU2D sub_56_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27655), 
          .S1(n898[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_1.INIT0 = 16'hF000;
    defparam sub_56_add_2_1.INIT1 = 16'h5555;
    defparam sub_56_add_2_1.INJECT1_0 = "NO";
    defparam sub_56_add_2_1.INJECT1_1 = "NO";
    LUT4 i24314_4_lut (.A(n11792), .B(count[9]), .C(n49_adj_122), .D(n30781), 
         .Z(n30668)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i24314_4_lut.init = 16'heeea;
    LUT4 i2_3_lut_adj_198 (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n49_adj_122)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_adj_198.init = 16'hfefe;
    LUT4 i24423_4_lut (.A(count[4]), .B(count[1]), .C(count[5]), .D(n30745), 
         .Z(n30781)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i24423_4_lut.init = 16'ha080;
    LUT4 i24387_3_lut (.A(count[0]), .B(count[2]), .C(count[3]), .Z(n30745)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24387_3_lut.init = 16'hfefe;
    LUT4 i24673_4_lut (.A(n30170), .B(n32497), .C(n32433), .D(n30548), 
         .Z(n30940)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i24673_4_lut.init = 16'h3031;
    LUT4 i2_4_lut (.A(n30761), .B(n32434), .C(n30347), .D(n30353), .Z(n30170)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;
    defparam i2_4_lut.init = 16'h5444;
    LUT4 i24403_3_lut (.A(n54), .B(n30668), .C(n23), .Z(n30761)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24403_3_lut.init = 16'hfefe;
    LUT4 i2_4_lut_adj_199 (.A(n30527), .B(count[9]), .C(n28414), .D(n4), 
         .Z(n30529)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_199.init = 16'hfeee;
    LUT4 i2_4_lut_adj_200 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28414)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_200.init = 16'hfeee;
    LUT4 i1_4_lut_rep_308 (.A(n11845), .B(count[13]), .C(count[12]), .D(n30529), 
         .Z(n32433)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_308.init = 16'heaaa;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n32457), .C(n30347), 
         .D(n30353), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i14448_2_lut (.A(n898[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14448_2_lut.init = 16'h8888;
    LUT4 i14447_2_lut (.A(n898[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14447_2_lut.init = 16'h8888;
    LUT4 i14446_2_lut (.A(n898[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14446_2_lut.init = 16'h8888;
    LUT4 i14445_2_lut (.A(n898[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14445_2_lut.init = 16'h8888;
    LUT4 i14444_2_lut (.A(n898[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14444_2_lut.init = 16'h8888;
    LUT4 i14443_2_lut (.A(n898[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14443_2_lut.init = 16'h8888;
    LUT4 i14442_2_lut (.A(n898[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14442_2_lut.init = 16'h8888;
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (n32378, n30431, databus, n224, 
            n3451, debug_c_c, register_addr, n30418, n32420, n3363, 
            n1318, n9, n1304, n1310, n12098, databus_out, \sendcount[1] , 
            \select[1] , n12788, n32472, n32395, n224_adj_42, n3181, 
            \select[2] , \select[4] , \select[7] , rw, \steps_reg[7] , 
            n9_adj_33, n4, debug_c_7, n32536, n11271, n5, n6, 
            \reg_size[2] , n32511, n34347, n32525, n30594, n11753, 
            \steps_reg[5] , n14, \steps_reg[3] , n15, \steps_reg[5]_adj_34 , 
            n14_adj_35, \steps_reg[3]_adj_36 , n15_adj_37, \steps_reg[5]_adj_38 , 
            n14_adj_39, \steps_reg[3]_adj_40 , n15_adj_41, debug_c_2, 
            debug_c_3, debug_c_4, debug_c_5, n34344, \reset_count[14] , 
            \reset_count[12] , \reset_count[13] , n30429, \reset_count[10] , 
            \reset_count[9] , n19896, n9395, GND_net, state, \rdata[0] , 
            n29195, \rdata[1] , n183, n32, bclk, n31583, n32436, 
            n32543, n32542, n32461, n9396_c, n31642) /* synthesis syn_module_defined=1 */ ;
    input n32378;
    input n30431;
    input [31:0]databus;
    input [31:0]n224;
    output [31:0]n3451;
    input debug_c_c;
    output [7:0]register_addr;
    input n30418;
    input n32420;
    output n3363;
    output n1318;
    output n9;
    output n1304;
    output n1310;
    input n12098;
    output [31:0]databus_out;
    output \sendcount[1] ;
    output \select[1] ;
    input n12788;
    output n32472;
    input n32395;
    input [31:0]n224_adj_42;
    output [31:0]n3181;
    output \select[2] ;
    output \select[4] ;
    output \select[7] ;
    output rw;
    input \steps_reg[7] ;
    output n9_adj_33;
    output n4;
    output debug_c_7;
    output n32536;
    input n11271;
    input n5;
    input n6;
    input \reg_size[2] ;
    input n32511;
    input n34347;
    input n32525;
    input n30594;
    output n11753;
    input \steps_reg[5] ;
    output n14;
    input \steps_reg[3] ;
    output n15;
    input \steps_reg[5]_adj_34 ;
    output n14_adj_35;
    input \steps_reg[3]_adj_36 ;
    output n15_adj_37;
    input \steps_reg[5]_adj_38 ;
    output n14_adj_39;
    input \steps_reg[3]_adj_40 ;
    output n15_adj_41;
    output debug_c_2;
    output debug_c_3;
    output debug_c_4;
    output debug_c_5;
    output n34344;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input \reset_count[13] ;
    input n30429;
    input \reset_count[10] ;
    input \reset_count[9] ;
    output n19896;
    output n9395;
    input GND_net;
    output [5:0]state;
    output \rdata[0] ;
    input n29195;
    output \rdata[1] ;
    input n183;
    output n32;
    output bclk;
    input n31583;
    input n32436;
    input n32543;
    input n32542;
    input n32461;
    input n9396_c;
    input n31642;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    
    wire n2497;
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    wire [31:0]n1286;
    wire [7:0]n2028;
    
    wire n8, n32535, n30, n30682;
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n32452, n32578, n33942, n14083;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n32450, n2539;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n14082;
    wire [3:0]n1682;
    
    wire n1687, n13423, n28418, n13424, n30300;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n30303, n29815, n32498, n11639, n30423, n29814;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n32440, n32415, n20305;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n11, n11_adj_10, n11_adj_11, n11_adj_12, n32474, n1391, 
        n11936;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n12022, n28273, n34346, n28268, n28280, n28265, n28283, 
        n29223, n29213, n29197, n29181, n29301, n29177, n29229, 
        n29231, n29179, n29297, n29299, n29303, n29355, n29225, 
        n29209, n30789, n30196, n11_adj_13, n11_adj_14, n11_adj_15, 
        n11_adj_16, n32545, n32546, n11_adj_17, n11_adj_18, n11_adj_19, 
        n11_adj_20, n10677, n9437, n29391, n10675, n9441, n1398, 
        n1397, n30136, n10751, n29441, n29501, n11_adj_21, n11_adj_22, 
        n32330, n2541, n11_adj_23, n11_adj_24, n32539, n32490, n4_c, 
        n32575;
    wire [7:0]n9241;
    
    wire n31647, n4_adj_25, n32571, n4_adj_26, n32565, n32505, n32439, 
        n5_c, n30199, n28369, n29211, n32552, n14425;
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n32551, n32555, n29818, n32554, n32558, n32557, n32561, 
        n32560, n32564, n32563, n32567, n32566, n32570, n32569, 
        n32574, n32573;
    wire [4:0]n18;
    wire [4:0]n19;
    
    wire n32577, n32576, n32507, n32562, n32328, n32329, n4_adj_30, 
        n32553, n4_adj_31, n32556, n4_adj_32, n32559, n4_adj_34, 
        n32568, n11539, n32494, n8679, escape, n9337, n30492, 
        n30493;
    wire [3:0]n8204;
    
    wire n14122, n32499, n30557, n32500, n32501, n9_adj_36, n32502, 
        n8_adj_38;
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n32324, n7, n32477, n30480, n30481, n32506, n28182, n17, 
        n9_adj_46, n31555, n31556, n32513, n32025, n32026, send, 
        n28397, n11238, n33939, n33940, n33941, n30202, n5_adj_56, 
        n30216, n28366, n14_c, n38, busy, n8_adj_60, n5_adj_62, 
        n30220, n28332, n18418, n6_c, n30201, n35, n30205, n55;
    wire [7:0]n4846;
    
    wire n30206, n30207, n5_adj_65, n30219, n28385, n7986, n28270, 
        n28279, n28258, n28351, n28333, n28227, n28253, n28324, 
        n28230, n28236, n28231, n28233, n28220, n28372, n28364, 
        n28371, n28398, n28213, n28342, n28313, n28367, n28330, 
        n28329, n1, n6_adj_66, n30208, n30775, n19966, n5_adj_71, 
        n30195, n30194, n30212, n30197, n30211, n30213, n30210, 
        n30209, n30200, n30214, n30769, n30215, n30217, n11477, 
        n6_adj_76, n30416, n30173, n6_adj_77, n5_adj_78, n30203, 
        n30221, n30222, n30223, n13_adj_80, n30225, n30218, n30224, 
        n30006, n5_adj_85, n30729, n5_adj_88, n5_adj_91, n30198, 
        n30131, n5_adj_92, n30204, n5_adj_93, n5_adj_94, n8_adj_95, 
        n4_adj_96, n6_adj_97, n6_adj_98, n15_adj_99, n30739, n5_adj_100, 
        n5_adj_101, n5_adj_102, n5_adj_103, n5_adj_104, n5_adj_105, 
        n29648, n5_adj_106, n5_adj_107, n5_adj_108, n5_adj_109, n5_adj_110, 
        n5_adj_111, n5_adj_112, n8_adj_113, n5_adj_114, n5_adj_115, 
        n5_adj_116, n5_adj_117, n5_adj_118, n5_adj_119, n5_adj_120;
    
    LUT4 mux_1384_i29_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[28]), 
         .D(n224[28]), .Z(n3451[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i28_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[27]), 
         .D(n224[27]), .Z(n3451[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_512_i5_3_lut (.A(n2497), .B(esc_data[4]), .C(n1286[18]), 
         .Z(n2028[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n1286[15]), .B(esc_data[7]), .C(n8), .D(esc_data[0]), 
         .Z(n2497)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'h2000;
    LUT4 i3_4_lut (.A(esc_data[2]), .B(n32535), .C(n30), .D(n30682), 
         .Z(n8)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut.init = 16'h3031;
    FD1S3IX bufcount__i3 (.D(n32578), .CK(debug_c_c), .CD(n32452), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_51 (.A(esc_data[1]), .B(esc_data[2]), .C(esc_data[4]), 
         .D(esc_data[3]), .Z(n30)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_51.init = 16'h2080;
    FD1S3IX bufcount__i2 (.D(n33942), .CK(debug_c_c), .CD(n32452), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n14083), .CK(debug_c_c), .CD(n32452), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2028[4]), .SP(n32450), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2028[3]), .SP(n32450), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2028[1]), .SP(n32450), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    LUT4 i24326_3_lut (.A(esc_data[1]), .B(esc_data[4]), .C(esc_data[3]), 
         .Z(n30682)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24326_3_lut.init = 16'hfefe;
    PFUMX i8317 (.BLUT(n14082), .ALUT(n1682[1]), .C0(n1687), .Z(n14083));
    PFUMX i7658 (.BLUT(n13423), .ALUT(n28418), .C0(n1687), .Z(n13424));
    LUT4 i2_4_lut (.A(n30300), .B(\buffer[0] [0]), .C(\buffer[0] [2]), 
         .D(\buffer[0] [1]), .Z(n30303)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'h8000;
    LUT4 mux_512_i4_3_lut (.A(n2497), .B(esc_data[3]), .C(n1286[18]), 
         .Z(n2028[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i4_3_lut.init = 16'hcaca;
    LUT4 mux_512_i2_3_lut (.A(n2497), .B(esc_data[1]), .C(n1286[18]), 
         .Z(n2028[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i2_3_lut.init = 16'hcaca;
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 mux_1384_i27_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[26]), 
         .D(n224[26]), .Z(n3451[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_4_lut (.A(\buffer[0] [0]), .B(n30300), .C(\buffer[0] [2]), 
         .D(\buffer[0] [1]), .Z(n29815)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32498), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n11639), .Z(n30423)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i2_3_lut_4_lut_adj_52 (.A(\buffer[0] [0]), .B(n30300), .C(\buffer[0] [1]), 
         .D(\buffer[0] [2]), .Z(n29814)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_52.init = 16'h0400;
    FD1P3IX sendcount__i0 (.D(n20305), .SP(n32440), .CD(n32415), .CK(debug_c_c), 
            .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_53 (.A(register_addr[4]), .B(register_addr[5]), .C(n30418), 
         .D(n32420), .Z(n3363)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_53.init = 16'h2000;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n32498), .C(\buffer[0] [7]), 
         .D(rx_data[7]), .Z(n11)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_54 (.A(bufcount[0]), .B(n32498), .C(\buffer[0] [6]), 
         .D(rx_data[6]), .Z(n11_adj_10)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_54.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_55 (.A(bufcount[0]), .B(n32498), .C(rx_data[5]), 
         .D(\buffer[0] [5]), .Z(n11_adj_11)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_55.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_56 (.A(bufcount[0]), .B(n32498), .C(rx_data[4]), 
         .D(\buffer[0] [4]), .Z(n11_adj_12)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_56.init = 16'hfe10;
    LUT4 reduce_or_453_i1_3_lut_4_lut (.A(n32474), .B(n11639), .C(\buffer[0] [7]), 
         .D(n1286[9]), .Z(n1391)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_453_i1_3_lut_4_lut.init = 16'hff80;
    FD1S3JX state_FSM_i1 (.D(n11936), .CK(debug_c_c), .PD(n32452), .Q(n1318));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n28273), .SP(n12022), .CD(n32452), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n28268), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n28280), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n28265), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n28283), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n29223), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n29213), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n29197), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n29181), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n29301), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n29177), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n29229), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n29231), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n29179), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n29297), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n29299), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n29303), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n29355), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n29225), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i2 (.D(n29209), .SP(n12022), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(n1286[3]), .B(n30789), .C(\buffer[2] [1]), 
         .Z(n30196)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i24_3_lut_4_lut_adj_57 (.A(bufcount[0]), .B(n32498), .C(rx_data[3]), 
         .D(\buffer[0] [3]), .Z(n11_adj_13)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_57.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_58 (.A(bufcount[0]), .B(n32498), .C(\buffer[0] [2]), 
         .D(rx_data[2]), .Z(n11_adj_14)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_58.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_59 (.A(bufcount[0]), .B(n32498), .C(\buffer[0] [1]), 
         .D(rx_data[1]), .Z(n11_adj_15)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_59.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_60 (.A(bufcount[0]), .B(n32498), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_adj_16)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_60.init = 16'hf1e0;
    PFUMX i25281 (.BLUT(n32545), .ALUT(n32546), .C0(sendcount[3]), .Z(n9));
    LUT4 i24_3_lut_4_lut_adj_61 (.A(bufcount[0]), .B(n32498), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_17)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_61.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_62 (.A(bufcount[0]), .B(n32498), .C(\buffer[1] [6]), 
         .D(rx_data[6]), .Z(n11_adj_18)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_62.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_63 (.A(bufcount[0]), .B(n32498), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_19)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_63.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_64 (.A(bufcount[0]), .B(n32498), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_20)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_64.init = 16'hf2d0;
    FD1S3IX state_FSM_i21 (.D(n10677), .CK(debug_c_c), .CD(n34346), .Q(n1286[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n9437), .CK(debug_c_c), .CD(n34346), .Q(n1286[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n29391), .CK(debug_c_c), .CD(n32452), .Q(n1286[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n10675), .CK(debug_c_c), .CD(n32452), .Q(n1286[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n9441), .CK(debug_c_c), .CD(n32452), .Q(n1286[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1398), .CK(debug_c_c), .CD(n32452), .Q(n1286[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1397), .CK(debug_c_c), .CD(n32452), .Q(n1304));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1286[12]), .CK(debug_c_c), .CD(n32452), 
            .Q(n1286[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1286[11]), .CK(debug_c_c), .CD(n32452), 
            .Q(n1286[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1286[10]), .CK(debug_c_c), .CD(n32452), 
            .Q(n1286[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1391), .CK(debug_c_c), .CD(n32452), .Q(n1286[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1310), .CK(debug_c_c), .CD(n32452), .Q(n1286[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1286[7]), .CK(debug_c_c), .CD(n32452), .Q(n1310));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1286[6]), .CK(debug_c_c), .CD(n32452), .Q(n1286[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1286[5]), .CK(debug_c_c), .CD(n32452), .Q(n1286[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n30423), .CK(debug_c_c), .CD(n32452), .Q(n1286[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n30136), .CK(debug_c_c), .CD(n32452), .Q(n1286[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n10751), .CK(debug_c_c), .CD(n32452), .Q(n1286[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n29441), .CK(debug_c_c), .CD(n32452), .Q(n1286[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i2 (.D(n29501), .CK(debug_c_c), .CD(n32452), .Q(n1286[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    LUT4 i24_3_lut_4_lut_adj_65 (.A(bufcount[0]), .B(n32498), .C(rx_data[3]), 
         .D(\buffer[1] [3]), .Z(n11_adj_21)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_65.init = 16'hfd20;
    FD1P3AX tx_data_i0_i0 (.D(n2028[0]), .SP(n32450), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n13424), .CK(debug_c_c), .CD(n32452), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    LUT4 i24_3_lut_4_lut_adj_66 (.A(bufcount[0]), .B(n32498), .C(\buffer[1] [2]), 
         .D(rx_data[2]), .Z(n11_adj_22)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_66.init = 16'hf2d0;
    FD1P3AX esc_data_i0_i0 (.D(n32330), .SP(n12098), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    LUT4 i24_3_lut_4_lut_adj_67 (.A(bufcount[0]), .B(n32498), .C(rx_data[1]), 
         .D(\buffer[1] [1]), .Z(n11_adj_23)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_67.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_68 (.A(bufcount[0]), .B(n32498), .C(rx_data[0]), 
         .D(\buffer[1] [0]), .Z(n11_adj_24)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_68.init = 16'hfd20;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n32539), .B(n32490), .C(n4_c), 
         .D(n32575), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 rx_data_3__bdd_4_lut_25823 (.A(rx_data[3]), .B(rx_data[2]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n31647)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_3__bdd_4_lut_25823.init = 16'h6001;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n32539), .B(n32490), .C(n4_adj_25), 
         .D(n32571), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n32539), .B(n32490), .C(n4_adj_26), 
         .D(n32565), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1286[4]), .B(n32505), .C(bufcount[0]), 
         .D(n32439), .Z(n28418)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hd222;
    LUT4 i2_4_lut_adj_69 (.A(databus[21]), .B(n5_c), .C(n1286[13]), .D(n30199), 
         .Z(n28369)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_69.init = 16'hffec;
    FD1P3IX buffer_0___i1 (.D(n29211), .SP(n12022), .CD(n32452), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 i24506_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n32552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24506_then_3_lut.init = 16'hcaca;
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    LUT4 i24506_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n32551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24506_else_3_lut.init = 16'hcaca;
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 i24509_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n32555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24509_then_3_lut.init = 16'hcaca;
    FD1P3AX select__i1 (.D(n29818), .SP(n12788), .CK(debug_c_c), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    LUT4 i24509_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n32554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24509_else_3_lut.init = 16'hcaca;
    LUT4 mux_1384_i17_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[16]), 
         .D(n224[16]), .Z(n3451[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i24512_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n32558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24512_then_3_lut.init = 16'hcaca;
    LUT4 i882_3_lut (.A(n1286[5]), .B(n32472), .C(n1286[10]), .Z(n2539)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i882_3_lut.init = 16'hc8c8;
    LUT4 mux_1314_i32_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[31]), 
         .D(n224_adj_42[31]), .Z(n3181[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 i24512_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n32557)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24512_else_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i31_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[30]), 
         .D(n224_adj_42[30]), .Z(n3181[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 i25248_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n32561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25248_then_3_lut.init = 16'hcaca;
    LUT4 i25248_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n32560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25248_else_3_lut.init = 16'hcaca;
    LUT4 i24515_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n32564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24515_then_3_lut.init = 16'hcaca;
    LUT4 i24515_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n32563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24515_else_3_lut.init = 16'hcaca;
    LUT4 i24518_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n32567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24518_then_3_lut.init = 16'hcaca;
    LUT4 i24518_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n32566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24518_else_3_lut.init = 16'hcaca;
    LUT4 i24521_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n32570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24521_then_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i30_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[29]), 
         .D(n224_adj_42[29]), .Z(n3181[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 i24521_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n32569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24521_else_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i29_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[28]), 
         .D(n224_adj_42[28]), .Z(n3181[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i28_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[27]), 
         .D(n224_adj_42[27]), .Z(n3181[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i28_3_lut_4_lut.init = 16'hf780;
    FD1P3AX select__i2 (.D(n29815), .SP(n12788), .CK(debug_c_c), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1P3AX select__i4 (.D(n29814), .SP(n12788), .CK(debug_c_c), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1P3AX select__i7 (.D(n30303), .SP(n12788), .CK(debug_c_c), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 i24524_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n32574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24524_then_3_lut.init = 16'hcaca;
    LUT4 i24524_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n32573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24524_else_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i27_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[26]), 
         .D(n224_adj_42[26]), .Z(n3181[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i27_3_lut_4_lut.init = 16'hf780;
    FD1P3AX sendcount__i2 (.D(n18[2]), .SP(n32440), .CK(debug_c_c), .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n19[1]), .SP(n32440), .CD(n32415), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 mux_1314_i26_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[25]), 
         .D(n224_adj_42[25]), .Z(n3181[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i25_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[24]), 
         .D(n224_adj_42[24]), .Z(n3181[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 i8325_then_4_lut (.A(bufcount[3]), .B(n1318), .C(n1286[3]), .D(n1286[4]), 
         .Z(n32577)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8325_then_4_lut.init = 16'haaa2;
    LUT4 i8325_else_4_lut (.A(bufcount[3]), .B(n1318), .C(n1286[3]), .D(n1286[4]), 
         .Z(n32576)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8325_else_4_lut.init = 16'h0002;
    LUT4 mux_1314_i24_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[23]), 
         .D(n224_adj_42[23]), .Z(n3181[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i23_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[22]), 
         .D(n224_adj_42[22]), .Z(n3181[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 n32328_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n32507), .C(n32562), 
         .D(n32328), .Z(n32329)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n32328_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 mux_1314_i22_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[21]), 
         .D(n224_adj_42[21]), .Z(n3181[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i21_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[20]), 
         .D(n224_adj_42[20]), .Z(n3181[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n32539), .B(n32490), .C(n4_adj_30), 
         .D(n32553), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n32539), .B(n32490), .C(n4_adj_31), 
         .D(n32556), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n32539), .B(n32490), .C(n4_adj_32), 
         .D(n32559), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_1314_i20_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[19]), 
         .D(n224_adj_42[19]), .Z(n3181[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i19_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[18]), 
         .D(n224_adj_42[18]), .Z(n3181[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i18_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[17]), 
         .D(n224_adj_42[17]), .Z(n3181[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i17_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[16]), 
         .D(n224_adj_42[16]), .Z(n3181[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i16_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[15]), 
         .D(n224_adj_42[15]), .Z(n3181[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n32539), .B(n32490), .C(n4_adj_34), 
         .D(n32568), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_1314_i15_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[14]), 
         .D(n224_adj_42[14]), .Z(n3181[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_70 (.A(rx_data[1]), .B(rx_data[4]), .C(rx_data[3]), 
         .Z(n11539)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_3_lut_adj_70.init = 16'h0808;
    LUT4 mux_1314_i14_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[13]), 
         .D(n224_adj_42[13]), .Z(n3181[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i13_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[12]), 
         .D(n224_adj_42[12]), .Z(n3181[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i14016_2_lut (.A(bufcount[1]), .B(n1318), .Z(n14082)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14016_2_lut.init = 16'h2222;
    LUT4 i2992_2_lut_rep_369 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32494)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2992_2_lut_rep_369.init = 16'h8888;
    FD1P3AX rw_498 (.D(n1286[10]), .SP(n2539), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i2891_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n8679)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2891_2_lut_3_lut.init = 16'h8080;
    FD1S3AX escape_501 (.D(n9337), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_71 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n30492)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_71.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_72 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n30493)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_72.init = 16'hbfbf;
    LUT4 mux_1314_i12_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[11]), 
         .D(n224_adj_42[11]), .Z(n3181[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i11_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[10]), 
         .D(n224_adj_42[10]), .Z(n3181[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i10_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[9]), 
         .D(n224_adj_42[9]), .Z(n3181[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i498_2_lut (.A(n1286[3]), .B(n1286[4]), .Z(n1687)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i498_2_lut.init = 16'heeee;
    LUT4 mux_1314_i9_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[8]), 
         .D(n224_adj_42[8]), .Z(n3181[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32546)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 mux_1384_i1_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[0]), 
         .D(n224[0]), .Z(n3451[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i8_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[7]), 
         .D(n224_adj_42[7]), .Z(n3181[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i16_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[15]), 
         .D(n224[15]), .Z(n3451[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i14794_3_lut_rep_325 (.A(n2497), .B(n32472), .C(n1286[18]), .Z(n32450)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i14794_3_lut_rep_325.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_73 (.A(n9), .B(n8204[0]), .C(n32472), .D(n1304), 
         .Z(n14425)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_73.init = 16'h8000;
    LUT4 i24678_2_lut_3_lut (.A(n2497), .B(n32472), .C(n1286[18]), .Z(n14122)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i24678_2_lut_3_lut.init = 16'h0808;
    LUT4 mux_1314_i7_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[6]), 
         .D(n224_adj_42[6]), .Z(n3181[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i6_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[5]), 
         .D(n224_adj_42[5]), .Z(n3181[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i2787_2_lut_rep_373 (.A(bufcount[1]), .B(bufcount[2]), .Z(n32498)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2787_2_lut_rep_373.init = 16'heeee;
    LUT4 i2424_2_lut_rep_349_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n32474)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2424_2_lut_rep_349_3_lut.init = 16'hfefe;
    LUT4 i4_2_lut_rep_374 (.A(n1304), .B(n1286[15]), .Z(n32499)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_374.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_74 (.A(n1304), .B(n1286[15]), .C(n1286[12]), 
         .Z(n30557)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_74.init = 16'hfefe;
    LUT4 i1_2_lut_rep_375 (.A(n1286[3]), .B(n1286[19]), .Z(n32500)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_375.init = 16'heeee;
    LUT4 mux_1314_i5_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[4]), 
         .D(n224_adj_42[4]), .Z(n3181[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_376 (.A(n1286[11]), .B(n1286[9]), .Z(n32501)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_376.init = 16'heeee;
    LUT4 i3_2_lut_3_lut_4_lut (.A(n1286[11]), .B(n1286[9]), .C(n1286[19]), 
         .D(n1286[3]), .Z(n9_adj_36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_512_i1_3_lut (.A(n2497), .B(esc_data[0]), .C(n1286[18]), 
         .Z(n2028[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i4_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[3]), 
         .D(n224_adj_42[3]), .Z(n3181[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i3_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[2]), 
         .D(n224_adj_42[2]), .Z(n3181[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut (.A(register_addr[1]), .B(\steps_reg[7] ), .Z(n9_adj_33)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_rep_377 (.A(n1286[13]), .B(n1286[7]), .C(n1286[5]), 
         .Z(n32502)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_rep_377.init = 16'hfefe;
    LUT4 i2_2_lut_4_lut (.A(n1286[13]), .B(n1286[7]), .C(n1286[5]), .D(n1286[17]), 
         .Z(n8_adj_38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut_4_lut.init = 16'hfffe;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_34)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 mux_1384_i15_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[14]), 
         .D(n224[14]), .Z(n3451[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i2_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[1]), 
         .D(n224_adj_42[1]), .Z(n3181[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i14_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[13]), 
         .D(n224[13]), .Z(n3451[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 n11281_bdd_2_lut (.A(sendcount[0]), .B(sendcount[3]), .Z(n32324)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n11281_bdd_2_lut.init = 16'hbbbb;
    LUT4 mux_1384_i13_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[12]), 
         .D(n224[12]), .Z(n3451[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i12_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[11]), 
         .D(n224[11]), .Z(n3451[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i11_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[10]), 
         .D(n224[10]), .Z(n3451[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i14686_3_lut_rep_380 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n32505)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i14686_3_lut_rep_380.init = 16'hecec;
    LUT4 mux_1384_i10_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[9]), 
         .D(n224[9]), .Z(n3451[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i9_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[8]), 
         .D(n224[8]), .Z(n3451[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_32)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1286[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hec00;
    LUT4 i2_2_lut_rep_352_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1286[4]), .Z(n32477)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_352_4_lut.init = 16'hecff;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_31)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_adj_75 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n30480)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_75.init = 16'hfbfb;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_30)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_adj_76 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n30481)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_76.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_381 (.A(n1304), .B(sendcount[4]), .Z(n32506)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_381.init = 16'h2222;
    FD1P3AX sendcount__i3 (.D(n28182), .SP(n32440), .CK(debug_c_c), .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3AX sendcount__i4 (.D(n17), .SP(n32440), .CK(debug_c_c), .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 i14458_4_lut (.A(sendcount[2]), .B(n32415), .C(n9_adj_46), .D(n32494), 
         .Z(n18[2])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14458_4_lut.init = 16'h1323;
    LUT4 expansion5_c_bdd_2_lut_24954_3_lut (.A(n1304), .B(sendcount[4]), 
         .C(n31555), .Z(n31556)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam expansion5_c_bdd_2_lut_24954_3_lut.init = 16'h2020;
    LUT4 mux_1384_i26_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[25]), 
         .D(n224[25]), .Z(n3451[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i25_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[24]), 
         .D(n224[24]), .Z(n3451[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_77 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_77.init = 16'h4444;
    LUT4 i13897_2_lut_rep_382 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32507)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13897_2_lut_rep_382.init = 16'heeee;
    LUT4 i1_2_lut_rep_365_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n32490)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_365_3_lut.init = 16'h1e1e;
    LUT4 mux_1384_i8_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[7]), 
         .D(n224[7]), .Z(n3451[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i7_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[6]), 
         .D(n224[6]), .Z(n3451[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i854_2_lut_rep_388 (.A(escape), .B(debug_c_7), .Z(n32513)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i854_2_lut_rep_388.init = 16'hbbbb;
    LUT4 i2_3_lut_rep_314_4_lut (.A(escape), .B(debug_c_7), .C(n30789), 
         .D(n1286[4]), .Z(n32439)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_314_4_lut.init = 16'hfffb;
    LUT4 i13895_2_lut (.A(sendcount[3]), .B(sendcount[0]), .Z(n8204[0])) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i13895_2_lut.init = 16'hdddd;
    LUT4 mux_1384_i6_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[5]), 
         .D(n224[5]), .Z(n3451[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i884_2_lut (.A(n1286[5]), .B(n32472), .Z(n2541)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i884_2_lut.init = 16'h8888;
    LUT4 mux_1384_i5_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[4]), 
         .D(n224[4]), .Z(n3451[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i4_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[3]), 
         .D(n224[3]), .Z(n3451[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 sendcount_4__bdd_3_lut_25127 (.A(sendcount[4]), .B(n32025), .C(sendcount[3]), 
         .Z(n32026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut_25127.init = 16'hcaca;
    LUT4 mux_1384_i20_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[19]), 
         .D(n224[19]), .Z(n3451[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 sendcount_4__bdd_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(sendcount[2]), 
         .D(\sendcount[1] ), .Z(n32025)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_4__bdd_4_lut.init = 16'h6aaa;
    FD1P3AX send_491 (.D(n11238), .SP(n28397), .CK(debug_c_c), .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 select_1742_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30492), .Z(n5_c)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 n30789_bdd_4_lut_25999 (.A(n30789), .B(n32513), .C(n1318), .D(n1286[3]), 
         .Z(n33939)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n30789_bdd_4_lut_25999.init = 16'hee0f;
    LUT4 n33939_bdd_2_lut (.A(n33939), .B(n1286[4]), .Z(n33940)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n33939_bdd_2_lut.init = 16'heeee;
    LUT4 n30789_bdd_4_lut (.A(bufcount[1]), .B(n1286[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n33941)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n30789_bdd_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_adj_78 (.A(n1286[3]), .B(n30789), .C(\buffer[2] [0]), 
         .Z(n30202)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_78.init = 16'h8080;
    LUT4 i2_4_lut_adj_79 (.A(databus[22]), .B(n5_adj_56), .C(n1286[13]), 
         .D(n30216), .Z(n28366)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_79.init = 16'hffec;
    LUT4 mux_1384_i3_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[2]), 
         .D(n224[2]), .Z(n3451[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i2_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[1]), 
         .D(n224[1]), .Z(n3451[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i32_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[31]), 
         .D(n224[31]), .Z(n3451[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i32_3_lut_4_lut.init = 16'hf780;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n32450), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_80 (.A(n1286[3]), .B(n30789), .C(n1286[13]), 
         .Z(n14_c)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_80.init = 16'hf8f8;
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n32450), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n32450), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_81 (.A(n38), .B(busy), .C(n31556), .D(n1286[17]), 
         .Z(n29391)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_81.init = 16'hfbfa;
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n32450), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 select_1742_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30492), .Z(n5_adj_56)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_82 (.A(n1286[15]), .B(esc_data[7]), .C(n8_adj_60), 
         .D(esc_data[0]), .Z(n38)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_82.init = 16'ha8aa;
    LUT4 mux_1384_i31_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[30]), 
         .D(n224[30]), .Z(n3451[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_83 (.A(databus[23]), .B(n5_adj_62), .C(n1286[13]), 
         .D(n30220), .Z(n28332)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_83.init = 16'hffec;
    LUT4 mux_1384_i30_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[29]), 
         .D(n224[29]), .Z(n3451[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_84 (.A(\buffer[0] [2]), .B(\buffer[0] [0]), .C(n30300), 
         .D(\buffer[0] [1]), .Z(n29818)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_4_lut_adj_84.init = 16'h0040;
    LUT4 i1_4_lut_adj_85 (.A(\buffer[0] [3]), .B(n18418), .C(n6_c), .D(\buffer[0] [4]), 
         .Z(n30300)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_85.init = 16'h0004;
    LUT4 i2_2_lut (.A(\buffer[0] [5]), .B(\buffer[0] [6]), .Z(n6_c)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_86 (.A(n1286[3]), .B(n30789), .C(\buffer[2] [5]), 
         .Z(n30201)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_86.init = 16'h8080;
    LUT4 i1_4_lut_adj_87 (.A(esc_data[1]), .B(esc_data[3]), .C(esc_data[4]), 
         .D(esc_data[2]), .Z(n35)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_87.init = 16'h5f4c;
    LUT4 i1_2_lut_3_lut_adj_88 (.A(n1286[3]), .B(n30789), .C(\buffer[2] [6]), 
         .Z(n30205)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_88.init = 16'h8080;
    LUT4 i51_4_lut (.A(esc_data[2]), .B(esc_data[3]), .C(esc_data[4]), 
         .D(esc_data[1]), .Z(n55)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i51_4_lut.init = 16'h9998;
    LUT4 i24332_2_lut_rep_410 (.A(esc_data[5]), .B(esc_data[6]), .Z(n32535)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24332_2_lut_rep_410.init = 16'heeee;
    LUT4 mux_1314_i1_3_lut_4_lut (.A(n32395), .B(n30418), .C(databus[0]), 
         .D(n224_adj_42[0]), .Z(n3181[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i3_3_lut_4_lut (.A(esc_data[5]), .B(esc_data[6]), .C(n55), .D(n35), 
         .Z(n8_adj_60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4912_3_lut (.A(busy), .B(n1286[17]), .C(n1286[16]), .Z(n10675)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4912_3_lut.init = 16'ha8a8;
    LUT4 select_1742_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30492), .Z(n5_adj_62)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_39_i5_4_lut.init = 16'h88c0;
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i4 (.D(n4846[4]), .SP(n12098), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n4846[2]), .SP(n12098), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n4846[1]), .SP(n12098), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_411 (.A(n1286[6]), .B(n1286[11]), .Z(n32536)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_411.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_89 (.A(n1286[6]), .B(n1286[11]), .C(n32472), 
         .Z(n18418)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_89.init = 16'he0e0;
    LUT4 i2882_2_lut_rep_414 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32539)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i2882_2_lut_rep_414.init = 16'h9999;
    LUT4 i1_2_lut_3_lut_adj_90 (.A(n1286[3]), .B(n30789), .C(\buffer[2] [7]), 
         .Z(n30206)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_90.init = 16'h8080;
    LUT4 i3680_3_lut (.A(n1286[16]), .B(n2497), .C(busy), .Z(n9441)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3680_3_lut.init = 16'hcece;
    LUT4 n11281_bdd_4_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(\buffer[5] [0]), 
         .D(\buffer[4] [0]), .Z(n32328)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n11281_bdd_4_lut_4_lut.init = 16'h6420;
    LUT4 i1_2_lut_3_lut_adj_91 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [0]), 
         .Z(n30207)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_91.init = 16'h8080;
    LUT4 i13896_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_adj_46), .Z(n19[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i13896_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 i2_4_lut_adj_92 (.A(databus[24]), .B(n5_adj_65), .C(n1286[13]), 
         .D(n30219), .Z(n28385)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_92.init = 16'hffec;
    FD1P3IX buffer_0___i22 (.D(n28270), .SP(n7986), .CD(n32452), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    LUT4 select_1742_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30493), .Z(n5_adj_65)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 i461_2_lut (.A(n9), .B(n1304), .Z(n1398)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i461_2_lut.init = 16'h4444;
    LUT4 i24686_2_lut (.A(sendcount[0]), .B(n9_adj_46), .Z(n20305)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24686_2_lut.init = 16'h7777;
    FD1P3IX buffer_0___i23 (.D(n28279), .SP(n7986), .CD(n32452), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n28258), .SP(n7986), .CD(n32452), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n28351), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n28333), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n28227), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n28253), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n28324), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n28230), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n28236), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n28231), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n28233), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n28220), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n28372), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n28364), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n28371), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n28369), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n28366), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n28332), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n28385), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n28398), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n28213), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n28342), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n28313), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n28367), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n28330), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n28329), .SP(n7986), .CD(n34346), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_93 (.A(sendcount[4]), .B(n1), .C(n6_adj_66), .D(n11271), 
         .Z(n9_adj_46)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_93.init = 16'hfeff;
    LUT4 equal_48_i1_3_lut (.A(sendcount[0]), .B(n5), .C(n6), .Z(n1)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_48_i1_3_lut.init = 16'h5656;
    LUT4 i1_2_lut_3_lut_adj_94 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [1]), 
         .Z(n30208)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_94.init = 16'h8080;
    LUT4 i2_4_lut_adj_95 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n32511), .Z(n6_adj_66)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_95.init = 16'he7de;
    LUT4 mux_1384_i24_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[23]), 
         .D(n224[23]), .Z(n3451[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i23_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[22]), 
         .D(n224[22]), .Z(n3451[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i23_3_lut_4_lut.init = 16'hf780;
    PFUMX i26000 (.BLUT(n33941), .ALUT(n33940), .C0(bufcount[2]), .Z(n33942));
    LUT4 i24431_4_lut (.A(rx_data[0]), .B(n30775), .C(rx_data[4]), .D(n19966), 
         .Z(n30789)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i24431_4_lut.init = 16'hfffd;
    LUT4 i2_4_lut_adj_96 (.A(databus[25]), .B(n5_adj_71), .C(n1286[13]), 
         .D(n30195), .Z(n28398)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_96.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_adj_97 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [2]), 
         .Z(n30194)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_97.init = 16'h8080;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32545)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 i1_2_lut_3_lut_adj_98 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [3]), 
         .Z(n30212)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_98.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_99 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [4]), 
         .Z(n30197)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_99.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_100 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [5]), 
         .Z(n30211)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_100.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_101 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [6]), 
         .Z(n30213)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_101.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_102 (.A(n1286[3]), .B(n30789), .C(\buffer[3] [7]), 
         .Z(n30210)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_102.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_103 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [0]), 
         .Z(n30209)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_103.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_104 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [1]), 
         .Z(n30200)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_104.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_105 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [2]), 
         .Z(n30214)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_105.init = 16'h8080;
    LUT4 mux_1384_i22_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[21]), 
         .D(n224[21]), .Z(n3451[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i21_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[20]), 
         .D(n224[20]), .Z(n3451[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 reduce_or_459_i1_3_lut (.A(busy), .B(n1286[13]), .C(n1286[20]), 
         .Z(n1397)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_459_i1_3_lut.init = 16'hdcdc;
    PFUMX i25250 (.BLUT(n32329), .ALUT(n32324), .C0(n9), .Z(n32330));
    LUT4 i24417_3_lut (.A(rx_data[3]), .B(n30769), .C(rx_data[1]), .Z(n30775)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24417_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_106 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [3]), 
         .Z(n30215)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_106.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_107 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [4]), 
         .Z(n30217)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_107.init = 16'h8080;
    LUT4 mux_1384_i19_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[18]), 
         .D(n224[18]), .Z(n3451[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_108 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [5]), 
         .Z(n30199)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_108.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_109 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [6]), 
         .Z(n30216)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_109.init = 16'h8080;
    LUT4 mux_1384_i18_3_lut_4_lut (.A(n32378), .B(n30431), .C(databus[17]), 
         .D(n224[17]), .Z(n3451[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i24411_3_lut (.A(rx_data[5]), .B(rx_data[7]), .C(rx_data[6]), 
         .Z(n30769)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24411_3_lut.init = 16'hfefe;
    LUT4 i7972_4_lut (.A(escape), .B(n11477), .C(n6_adj_76), .D(n1286[3]), 
         .Z(n9337)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i7972_4_lut.init = 16'h1aaa;
    LUT4 i1_2_lut_3_lut_adj_110 (.A(n1286[3]), .B(n30789), .C(\buffer[4] [7]), 
         .Z(n30220)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_110.init = 16'h8080;
    LUT4 i2_2_lut_adj_111 (.A(debug_c_7), .B(n32472), .Z(n6_adj_76)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_111.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_112 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [0]), 
         .Z(n30219)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_112.init = 16'h8080;
    LUT4 i14237_2_lut (.A(rx_data[2]), .B(rx_data[1]), .Z(n19966)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14237_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_113 (.A(n30416), .B(debug_c_7), .C(n1318), .D(n1286[1]), 
         .Z(n11936)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_113.init = 16'hbbba;
    LUT4 i3_4_lut_adj_114 (.A(n34347), .B(n32525), .C(register_addr[2]), 
         .D(n30594), .Z(n11753)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_adj_114.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_adj_115 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [1]), 
         .Z(n30195)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_115.init = 16'h8080;
    LUT4 i4_4_lut (.A(rx_data[2]), .B(n30173), .C(rx_data[5]), .D(n6_adj_77), 
         .Z(n11639)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i4_4_lut.init = 16'h0800;
    LUT4 i3_4_lut_adj_116 (.A(sendcount[3]), .B(n32507), .C(sendcount[2]), 
         .D(n32506), .Z(n30416)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_116.init = 16'h0200;
    LUT4 select_1742_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30493), .Z(n5_adj_71)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_117 (.A(databus[4]), .B(n5_adj_78), .C(n1286[13]), 
         .D(n30203), .Z(n28273)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_117.init = 16'hffec;
    LUT4 i1_2_lut_adj_118 (.A(register_addr[1]), .B(\steps_reg[5] ), .Z(n14)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_118.init = 16'h8888;
    LUT4 select_1742_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30480), .Z(n5_adj_78)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_119 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [2]), 
         .Z(n30221)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_119.init = 16'h8080;
    LUT4 i1_2_lut_adj_120 (.A(register_addr[1]), .B(\steps_reg[3] ), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_120.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_121 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [3]), 
         .Z(n30222)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_121.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_122 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [4]), 
         .Z(n30223)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_122.init = 16'h8080;
    LUT4 i2_4_lut_adj_123 (.A(escape), .B(n13_adj_80), .C(debug_c_7), 
         .D(n11539), .Z(n30173)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2_4_lut_adj_123.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_124 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [5]), 
         .Z(n30225)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_124.init = 16'h8080;
    LUT4 i1_2_lut_adj_125 (.A(n1286[3]), .B(rx_data[0]), .Z(n6_adj_77)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_adj_125.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_126 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [6]), 
         .Z(n30218)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_126.init = 16'h8080;
    LUT4 i1_2_lut_adj_127 (.A(register_addr[1]), .B(\steps_reg[5]_adj_34 ), 
         .Z(n14_adj_35)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_127.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_128 (.A(n1286[3]), .B(n30789), .C(\buffer[5] [7]), 
         .Z(n30224)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_128.init = 16'h8080;
    LUT4 i1_2_lut_adj_129 (.A(register_addr[1]), .B(\steps_reg[3]_adj_36 ), 
         .Z(n15_adj_37)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_129.init = 16'h8888;
    LUT4 i2_4_lut_adj_130 (.A(n32415), .B(sendcount[3]), .C(n9_adj_46), 
         .D(n8679), .Z(n28182)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_130.init = 16'h1040;
    LUT4 equal_143_i13_2_lut (.A(rx_data[6]), .B(rx_data[7]), .Z(n13_adj_80)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam equal_143_i13_2_lut.init = 16'heeee;
    LUT4 i13991_2_lut (.A(bufcount[0]), .B(n1318), .Z(n13423)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i13991_2_lut.init = 16'h2222;
    LUT4 i24810_3_lut (.A(debug_c_7), .B(n30006), .C(n1286[3]), .Z(n30136)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i24810_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_adj_131 (.A(n1286[4]), .B(\buffer[0] [0]), .C(n11_adj_16), 
         .D(n14_c), .Z(n29211)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_131.init = 16'heca0;
    LUT4 i2_4_lut_adj_132 (.A(databus[26]), .B(n5_adj_85), .C(n1286[13]), 
         .D(n30221), .Z(n28213)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_132.init = 16'hffec;
    LUT4 select_1742_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30493), .Z(n5_adj_85)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 i24765_2_lut_2_lut (.A(n32472), .B(n7986), .Z(n12022)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i24765_2_lut_2_lut.init = 16'hdddd;
    LUT4 i24801_4_lut (.A(n7), .B(n30729), .C(n32513), .D(n1286[3]), 
         .Z(n7986)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i24801_4_lut.init = 16'h0544;
    LUT4 i1_2_lut_adj_133 (.A(register_addr[1]), .B(\steps_reg[5]_adj_38 ), 
         .Z(n14_adj_39)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_133.init = 16'h8888;
    LUT4 i2_4_lut_adj_134 (.A(databus[27]), .B(n5_adj_88), .C(n1286[13]), 
         .D(n30222), .Z(n28342)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_134.init = 16'hffec;
    LUT4 i3_4_lut_adj_135 (.A(n30769), .B(n31647), .C(rx_data[0]), .D(escape), 
         .Z(n30006)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_135.init = 16'h0040;
    LUT4 i24371_3_lut (.A(n1286[13]), .B(n1318), .C(n1286[4]), .Z(n30729)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24371_3_lut.init = 16'hfefe;
    LUT4 select_1742_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30493), .Z(n5_adj_88)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_adj_136 (.A(register_addr[1]), .B(\steps_reg[3]_adj_40 ), 
         .Z(n15_adj_41)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_136.init = 16'h8888;
    LUT4 i2_4_lut_adj_137 (.A(databus[3]), .B(n5_adj_91), .C(n1286[13]), 
         .D(n30198), .Z(n28268)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_137.init = 16'hffec;
    LUT4 i4986_3_lut (.A(debug_c_7), .B(n1286[3]), .C(n1286[2]), .Z(n10751)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4986_3_lut.init = 16'h5454;
    LUT4 select_1742_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30480), .Z(n5_adj_91)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_138 (.A(n1286[4]), .B(debug_c_7), .C(n1286[2]), 
         .D(n30131), .Z(n29441)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_138.init = 16'heeea;
    LUT4 i2_4_lut_adj_139 (.A(databus[2]), .B(n5_adj_92), .C(n1286[13]), 
         .D(n30204), .Z(n28280)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_139.init = 16'hffec;
    LUT4 select_1742_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30480), .Z(n5_adj_92)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_140 (.A(databus[1]), .B(n5_adj_93), .C(n1286[13]), 
         .D(n30196), .Z(n28265)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_140.init = 16'hffec;
    LUT4 select_1742_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30480), .Z(n5_adj_93)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i2_3_lut (.A(n1286[19]), .B(n1286[16]), .C(n11238), .Z(n28397)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i2_3_lut.init = 16'hefef;
    LUT4 i24808_3_lut (.A(n32472), .B(n1286[20]), .C(n1286[17]), .Z(n11238)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i24808_3_lut.init = 16'h0202;
    LUT4 mux_1578_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n9), .Z(n4846[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1578_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_26)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 mux_1578_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n9), .Z(n4846[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1578_i3_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_141 (.A(databus[0]), .B(n5_adj_94), .C(n1286[13]), 
         .D(n30202), .Z(n28283)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_141.init = 16'hffec;
    LUT4 select_1742_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30480), .Z(n5_adj_94)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_25)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 mux_1578_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n9), .Z(n4846[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1578_i2_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_c)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 i5_4_lut (.A(n9_adj_36), .B(n1286[15]), .C(n8_adj_38), .D(n1286[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_142 (.A(n1286[2]), .B(n32499), .C(n8_adj_95), .D(n1286[18]), 
         .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_142.init = 16'hfffe;
    LUT4 i3_4_lut_adj_143 (.A(n32500), .B(n1286[10]), .C(n4_adj_96), .D(n1286[6]), 
         .Z(n8_adj_95)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_143.init = 16'hfffe;
    LUT4 i1_2_lut_adj_144 (.A(n1286[11]), .B(n1286[7]), .Z(n4_adj_96)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_144.init = 16'heeee;
    LUT4 i4_4_lut_adj_145 (.A(n1286[20]), .B(n30557), .C(n32502), .D(n6_adj_97), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4_4_lut_adj_145.init = 16'hfffe;
    LUT4 i1_2_lut_adj_146 (.A(n1286[4]), .B(n1286[6]), .Z(n6_adj_97)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_146.init = 16'heeee;
    LUT4 i4_4_lut_adj_147 (.A(n1310), .B(n30557), .C(n32501), .D(n6_adj_98), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_147.init = 16'hfffe;
    LUT4 i1_4_lut_adj_148 (.A(n15_adj_99), .B(n1286[3]), .C(n1318), .D(n30739), 
         .Z(n30131)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_148.init = 16'h50dc;
    LUT4 i1_2_lut_adj_149 (.A(n1286[13]), .B(n1286[10]), .Z(n6_adj_98)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_149.init = 16'heeee;
    LUT4 i2_4_lut_adj_150 (.A(databus[28]), .B(n5_adj_100), .C(n1286[13]), 
         .D(n30223), .Z(n28313)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_150.init = 16'hffec;
    LUT4 i1_4_lut_adj_151 (.A(n1286[4]), .B(\buffer[1] [7]), .C(n11_adj_17), 
         .D(n14_c), .Z(n29223)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_151.init = 16'heca0;
    LUT4 select_1742_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30493), .Z(n5_adj_100)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_152 (.A(n1286[4]), .B(\buffer[1] [6]), .C(n11_adj_18), 
         .D(n14_c), .Z(n29213)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_152.init = 16'heca0;
    LUT4 i2_4_lut_adj_153 (.A(databus[29]), .B(n5_adj_101), .C(n1286[13]), 
         .D(n30225), .Z(n28367)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_153.init = 16'hffec;
    LUT4 i1_4_lut_adj_154 (.A(n1286[4]), .B(\buffer[1] [5]), .C(n11_adj_19), 
         .D(n14_c), .Z(n29197)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_154.init = 16'heca0;
    LUT4 i2_4_lut_adj_155 (.A(databus[5]), .B(n5_adj_102), .C(n1286[13]), 
         .D(n30201), .Z(n28270)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_155.init = 16'hffec;
    LUT4 select_1742_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30480), .Z(n5_adj_102)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_156 (.A(databus[6]), .B(n5_adj_103), .C(n1286[13]), 
         .D(n30205), .Z(n28279)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_156.init = 16'hffec;
    LUT4 select_1742_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30480), .Z(n5_adj_103)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 select_1742_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30493), .Z(n5_adj_101)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_157 (.A(n1286[4]), .B(\buffer[1] [4]), .C(n11_adj_20), 
         .D(n14_c), .Z(n29181)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_157.init = 16'heca0;
    LUT4 i2_4_lut_adj_158 (.A(databus[7]), .B(n5_adj_104), .C(n1286[13]), 
         .D(n30206), .Z(n28258)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_158.init = 16'hffec;
    LUT4 select_1742_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30480), .Z(n5_adj_104)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_159 (.A(databus[8]), .B(n5_adj_105), .C(n1286[13]), 
         .D(n30207), .Z(n28351)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_159.init = 16'hffec;
    LUT4 select_1742_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30481), .Z(n5_adj_105)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 i24381_3_lut (.A(n11477), .B(escape), .C(n15_adj_99), .Z(n30739)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24381_3_lut.init = 16'hecec;
    LUT4 n30415_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n31555)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n30415_bdd_4_lut.init = 16'h4001;
    LUT4 i1_4_lut_adj_160 (.A(n1286[4]), .B(\buffer[1] [3]), .C(n11_adj_21), 
         .D(n14_c), .Z(n29301)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_160.init = 16'heca0;
    LUT4 i2_4_lut_adj_161 (.A(n29648), .B(rx_data[4]), .C(rx_data[1]), 
         .D(rx_data[3]), .Z(n11477)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(150[12:17])
    defparam i2_4_lut_adj_161.init = 16'hbfff;
    LUT4 i2_4_lut_adj_162 (.A(databus[9]), .B(n5_adj_106), .C(n1286[13]), 
         .D(n30208), .Z(n28333)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_162.init = 16'hffec;
    LUT4 select_1742_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30481), .Z(n5_adj_106)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_163 (.A(n1286[4]), .B(\buffer[1] [2]), .C(n11_adj_22), 
         .D(n14_c), .Z(n29177)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_163.init = 16'heca0;
    LUT4 i2_4_lut_adj_164 (.A(databus[10]), .B(n5_adj_107), .C(n1286[13]), 
         .D(n30194), .Z(n28227)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_164.init = 16'hffec;
    LUT4 select_1742_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30481), .Z(n5_adj_107)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_165 (.A(n1286[4]), .B(\buffer[1] [1]), .C(n11_adj_23), 
         .D(n14_c), .Z(n29229)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_165.init = 16'heca0;
    LUT4 i2_4_lut_adj_166 (.A(databus[30]), .B(n5_adj_108), .C(n1286[13]), 
         .D(n30218), .Z(n28330)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_166.init = 16'hffec;
    LUT4 i2_4_lut_adj_167 (.A(databus[11]), .B(n5_adj_109), .C(n1286[13]), 
         .D(n30212), .Z(n28253)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_167.init = 16'hffec;
    LUT4 select_1742_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30481), .Z(n5_adj_109)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i3_4_lut_adj_168 (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), 
         .D(n29648), .Z(n15_adj_99)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(150[12:17])
    defparam i3_4_lut_adj_168.init = 16'hfffe;
    LUT4 i2_4_lut_adj_169 (.A(n13_adj_80), .B(rx_data[5]), .C(rx_data[2]), 
         .D(rx_data[0]), .Z(n29648)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(150[12:17])
    defparam i2_4_lut_adj_169.init = 16'hfeff;
    LUT4 i1_4_lut_adj_170 (.A(n1286[4]), .B(\buffer[1] [0]), .C(n11_adj_24), 
         .D(n14_c), .Z(n29231)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_170.init = 16'heca0;
    LUT4 select_1742_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30493), .Z(n5_adj_108)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_171 (.A(databus[12]), .B(n5_adj_110), .C(n1286[13]), 
         .D(n30197), .Z(n28324)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_171.init = 16'hffec;
    LUT4 i1_4_lut_adj_172 (.A(n1286[4]), .B(\buffer[0] [7]), .C(n11), 
         .D(n14_c), .Z(n29179)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_172.init = 16'heca0;
    LUT4 select_1742_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30481), .Z(n5_adj_110)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_173 (.A(databus[31]), .B(n5_adj_111), .C(n1286[13]), 
         .D(n30224), .Z(n28329)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_173.init = 16'hffec;
    LUT4 i1_4_lut_adj_174 (.A(n1286[4]), .B(\buffer[0] [6]), .C(n11_adj_10), 
         .D(n14_c), .Z(n29297)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_174.init = 16'heca0;
    LUT4 i2_4_lut_adj_175 (.A(databus[13]), .B(n5_adj_112), .C(n1286[13]), 
         .D(n30211), .Z(n28230)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_175.init = 16'hffec;
    LUT4 i1_4_lut_adj_176 (.A(n1286[4]), .B(\buffer[0] [5]), .C(n11_adj_11), 
         .D(n14_c), .Z(n29299)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_176.init = 16'heca0;
    LUT4 select_1742_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30481), .Z(n5_adj_112)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 select_1742_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30493), .Z(n5_adj_111)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_177 (.A(n32474), .B(debug_c_7), .C(n11639), .D(n8_adj_113), 
         .Z(n29501)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_177.init = 16'hdc50;
    LUT4 i2_4_lut_adj_178 (.A(databus[14]), .B(n5_adj_114), .C(n1286[13]), 
         .D(n30213), .Z(n28236)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_178.init = 16'hffec;
    LUT4 i1_3_lut (.A(n15_adj_99), .B(n1286[1]), .C(n1318), .Z(n8_adj_113)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 select_1742_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30481), .Z(n5_adj_114)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_179 (.A(databus[15]), .B(n5_adj_115), .C(n1286[13]), 
         .D(n30210), .Z(n28231)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_179.init = 16'hffec;
    LUT4 select_1742_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30481), .Z(n5_adj_115)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i4913_3_lut (.A(busy), .B(n1286[20]), .C(n1286[19]), .Z(n10677)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4913_3_lut.init = 16'ha8a8;
    LUT4 i14792_3_lut_rep_315 (.A(n1286[13]), .B(n32472), .C(n1304), .Z(n32440)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i14792_3_lut_rep_315.init = 16'hc8c8;
    LUT4 i2_4_lut_adj_180 (.A(databus[16]), .B(n5_adj_116), .C(n1286[13]), 
         .D(n30209), .Z(n28233)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_180.init = 16'hffec;
    LUT4 select_1742_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30492), .Z(n5_adj_116)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_181 (.A(n1286[4]), .B(\buffer[0] [4]), .C(n11_adj_12), 
         .D(n14_c), .Z(n29303)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_181.init = 16'heca0;
    LUT4 i2_4_lut_adj_182 (.A(databus[17]), .B(n5_adj_117), .C(n1286[13]), 
         .D(n30200), .Z(n28220)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_182.init = 16'hffec;
    LUT4 i24779_2_lut_3_lut_4_lut (.A(n1286[13]), .B(n32472), .C(n1304), 
         .D(n32026), .Z(n17)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i24779_2_lut_3_lut_4_lut.init = 16'hf700;
    LUT4 i1_4_lut_adj_183 (.A(n1286[4]), .B(\buffer[0] [3]), .C(n11_adj_13), 
         .D(n14_c), .Z(n29355)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_183.init = 16'heca0;
    LUT4 i24690_2_lut_rep_290_3_lut (.A(n1286[13]), .B(n32472), .C(n1304), 
         .Z(n32415)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i24690_2_lut_rep_290_3_lut.init = 16'h0808;
    LUT4 i3676_3_lut (.A(n1286[19]), .B(n1286[18]), .C(busy), .Z(n9437)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3676_3_lut.init = 16'hcece;
    LUT4 select_1742_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30492), .Z(n5_adj_117)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_184 (.A(n1286[3]), .B(n30789), .C(\buffer[2] [4]), 
         .Z(n30203)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_184.init = 16'h8080;
    LUT4 i2_4_lut_adj_185 (.A(databus[18]), .B(n5_adj_118), .C(n1286[13]), 
         .D(n30214), .Z(n28372)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_185.init = 16'hffec;
    LUT4 select_1742_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30492), .Z(n5_adj_118)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_186 (.A(n1286[3]), .B(n30789), .C(\buffer[2] [3]), 
         .Z(n30198)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_186.init = 16'h8080;
    FD1P3AX rw_498_rep_420 (.D(n1286[10]), .SP(n2539), .CK(debug_c_c), 
            .Q(n34344));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_420.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_187 (.A(databus[19]), .B(n5_adj_119), .C(n1286[13]), 
         .D(n30215), .Z(n28364)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_187.init = 16'hffec;
    LUT4 select_1742_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30492), .Z(n5_adj_119)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_188 (.A(n1286[3]), .B(n30789), .C(\buffer[2] [2]), 
         .Z(n30204)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_188.init = 16'h8080;
    LUT4 i1_4_lut_adj_189 (.A(n1286[4]), .B(\buffer[0] [2]), .C(n11_adj_14), 
         .D(n14_c), .Z(n29225)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_189.init = 16'heca0;
    LUT4 i2_4_lut_adj_190 (.A(databus[20]), .B(n5_adj_120), .C(n1286[13]), 
         .D(n30217), .Z(n28371)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_190.init = 16'hffec;
    PFUMX i25301 (.BLUT(n32576), .ALUT(n32577), .C0(n32439), .Z(n32578));
    LUT4 i1_4_lut_adj_191 (.A(n1286[4]), .B(\buffer[0] [1]), .C(n11_adj_15), 
         .D(n14_c), .Z(n29209)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_191.init = 16'heca0;
    PFUMX i25299 (.BLUT(n32573), .ALUT(n32574), .C0(sendcount[0]), .Z(n32575));
    LUT4 select_1742_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30492), .Z(n5_adj_120)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_36_i5_4_lut.init = 16'h88c0;
    PFUMX i25297 (.BLUT(n32569), .ALUT(n32570), .C0(sendcount[0]), .Z(n32571));
    PFUMX i25295 (.BLUT(n32566), .ALUT(n32567), .C0(sendcount[0]), .Z(n32568));
    PFUMX i25293 (.BLUT(n32563), .ALUT(n32564), .C0(sendcount[0]), .Z(n32565));
    PFUMX i25291 (.BLUT(n32560), .ALUT(n32561), .C0(sendcount[0]), .Z(n32562));
    PFUMX i25289 (.BLUT(n32557), .ALUT(n32558), .C0(sendcount[0]), .Z(n32559));
    PFUMX i25287 (.BLUT(n32554), .ALUT(n32555), .C0(sendcount[0]), .Z(n32556));
    PFUMX i25285 (.BLUT(n32551), .ALUT(n32552), .C0(sendcount[0]), .Z(n32553));
    LUT4 i2838_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n32439), .C(n32477), 
         .D(bufcount[0]), .Z(n1682[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2838_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    \UARTTransmitter(baud_div=12)  uart_output (.\reset_count[14] (\reset_count[14] ), 
            .\reset_count[12] (\reset_count[12] ), .\reset_count[13] (\reset_count[13] ), 
            .n30429(n30429), .n32472(n32472), .n32452(n32452), .tx_data({tx_data}), 
            .send(send), .n34346(n34346), .busy(busy), .\reset_count[10] (\reset_count[10] ), 
            .\reset_count[9] (\reset_count[9] ), .n19896(n19896), .n9395(n9395), 
            .debug_c_c(debug_c_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.state({state}), .rdata({Open_46, 
            Open_47, Open_48, Open_49, Open_50, Open_51, Open_52, 
            \rdata[0] }), .debug_c_c(debug_c_c), .n32472(n32472), .rx_data({rx_data}), 
            .n32452(n32452), .n34346(n34346), .n29195(n29195), .\rdata[1] (\rdata[1] ), 
            .n183(n183), .n32(n32), .bclk(bclk), .debug_c_7(debug_c_7), 
            .n31583(n31583), .n32436(n32436), .n32543(n32543), .n32542(n32542), 
            .n32461(n32461), .n9396_c(n9396_c), .n31642(n31642), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (\reset_count[14] , \reset_count[12] , 
            \reset_count[13] , n30429, n32472, n32452, tx_data, send, 
            n34346, busy, \reset_count[10] , \reset_count[9] , n19896, 
            n9395, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input \reset_count[13] ;
    input n30429;
    output n32472;
    output n32452;
    input [7:0]tx_data;
    input send;
    output n34346;
    output busy;
    input \reset_count[10] ;
    input \reset_count[9] ;
    output n19896;
    output n9395;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n2, n30861;
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n7;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n10, n31581, n7984, n12208, n29073, n17, n17_adj_9, n104, 
        n31579, n31989, n31990, n13675, n30859, n30860, n31580, 
        n2533, n30391, n30390, n30246, n19773, n32428;
    
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n30861), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i14281_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i14281_4_lut.init = 16'hfcee;
    LUT4 i1_4_lut_rep_347 (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n30429), .Z(n32472)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_rep_347.init = 16'hfaea;
    LUT4 i14769_1_lut_rep_327_4_lut (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n30429), .Z(n32452)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;
    defparam i14769_1_lut_rep_327_4_lut.init = 16'h0515;
    FD1S3IX state__i0 (.D(n31581), .CK(bclk), .CD(n32452), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n7984), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n7984), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n7984), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n7984), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n7984), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n7984), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n7984), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n7984), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX state__i3 (.D(n29073), .SP(n12208), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 i24_4_lut_4_lut (.A(state[3]), .B(state[0]), .C(state[1]), .D(send), 
         .Z(n17_adj_9)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i24_4_lut_4_lut.init = 16'h8001;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    LUT4 state_1__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n31579)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 i14769_1_lut_rep_422 (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n30429), .Z(n34346)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;
    defparam i14769_1_lut_rep_422.init = 16'h0515;
    LUT4 state_2__bdd_4_lut_25115 (.A(state[0]), .B(state[3]), .C(state[1]), 
         .D(send), .Z(n31989)) /* synthesis lut_function=(A (B (C))+!A !(B+(C+!(D)))) */ ;
    defparam state_2__bdd_4_lut_25115.init = 16'h8180;
    LUT4 n31989_bdd_2_lut (.A(n31989), .B(state[2]), .Z(n31990)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n31989_bdd_2_lut.init = 16'h2222;
    FD1P3IX busy_34 (.D(n13675), .SP(n31990), .CD(n34346), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    PFUMX i24503 (.BLUT(n30859), .ALUT(n30860), .C0(state[1]), .Z(n30861));
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(send), .Z(n31580)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8f0e;
    LUT4 i1_2_lut (.A(state[0]), .B(state[1]), .Z(n2533)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_49 (.A(\reset_count[10] ), .B(\reset_count[9] ), .Z(n19896)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_49.init = 16'h8888;
    FD1P3AX state__i1 (.D(n30391), .SP(n12208), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX state__i2 (.D(n30390), .SP(n12208), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n32452), .CK(bclk), .Q(n9395)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n30246), .B(state[2]), .C(n19773), .D(n32472), 
         .Z(n7984)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_adj_50 (.A(send), .B(state[3]), .Z(n30246)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_50.init = 16'h2222;
    LUT4 i14044_2_lut (.A(state[1]), .B(state[0]), .Z(n19773)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14044_2_lut.init = 16'heeee;
    LUT4 i24816_3_lut (.A(n32472), .B(n17_adj_9), .C(state[2]), .Z(n12208)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i24816_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut (.A(n32472), .B(state[3]), .C(state[2]), .D(n2533), 
         .Z(n29073)) /* synthesis lut_function=(!((B (C)+!B !(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h2808;
    LUT4 i8330_1_lut (.A(state[3]), .Z(n13675)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i8330_1_lut.init = 16'h5555;
    LUT4 i24501_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n30859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24501_3_lut.init = 16'hcaca;
    LUT4 i24502_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n30860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24502_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_303 (.A(n32472), .B(state[2]), .C(state[3]), .Z(n32428)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut_rep_303.init = 16'h2a2a;
    LUT4 i1_3_lut_4_lut (.A(n32472), .B(state[2]), .C(state[3]), .D(n2533), 
         .Z(n30390)) /* synthesis lut_function=(!((B (C+(D))+!B !(D))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2208;
    PFUMX i24955 (.BLUT(n31580), .ALUT(n31579), .C0(state[2]), .Z(n31581));
    LUT4 i1_3_lut (.A(state[1]), .B(n32428), .C(state[0]), .Z(n30391)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    \ClockDividerP(factor=12)  baud_gen (.debug_c_c(debug_c_c), .bclk(bclk), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (debug_c_c, bclk, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output bclk;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    
    wire n55;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n56, n4, n14394, n52, n44, n35, n54, n48, n36, n46, 
        n32, n50, n40;
    wire [31:0]n102;
    
    wire n7264, n27535, n27536, n27922, n27921, n27920, n27919, 
        n27918, n27917, n27916, n27915, n27914, n27913, n27912, 
        n27911, n27910, n27909, n27908, n27907, n27550, n27549, 
        n27548, n27547, n27546, n27545, n27544, n27543, n27542, 
        n27541, n27540, n27539, n27538, n27537;
    
    LUT4 i24789_4_lut (.A(n55), .B(count[1]), .C(n56), .D(n4), .Z(n14394)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24789_4_lut.init = 16'h0400;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[3]), .B(count[0]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i11_2_lut.init = 16'heeee;
    FD1S3IX count_2181__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i0.GSR = "ENABLED";
    FD1S3AX clk_o_14 (.D(n7264), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D sub_1736_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27535), .COUT(n27536));
    defparam sub_1736_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1736_add_2_4.INIT1 = 16'h5555;
    defparam sub_1736_add_2_4.INJECT1_0 = "NO";
    defparam sub_1736_add_2_4.INJECT1_1 = "NO";
    FD1S3IX count_2181__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i1.GSR = "ENABLED";
    FD1S3IX count_2181__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i2.GSR = "ENABLED";
    FD1S3IX count_2181__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i3.GSR = "ENABLED";
    FD1S3IX count_2181__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i4.GSR = "ENABLED";
    FD1S3IX count_2181__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i5.GSR = "ENABLED";
    FD1S3IX count_2181__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i6.GSR = "ENABLED";
    FD1S3IX count_2181__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i7.GSR = "ENABLED";
    FD1S3IX count_2181__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i8.GSR = "ENABLED";
    FD1S3IX count_2181__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i9.GSR = "ENABLED";
    FD1S3IX count_2181__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i10.GSR = "ENABLED";
    FD1S3IX count_2181__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i11.GSR = "ENABLED";
    FD1S3IX count_2181__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i12.GSR = "ENABLED";
    FD1S3IX count_2181__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i13.GSR = "ENABLED";
    FD1S3IX count_2181__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i14.GSR = "ENABLED";
    FD1S3IX count_2181__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i15.GSR = "ENABLED";
    FD1S3IX count_2181__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i16.GSR = "ENABLED";
    FD1S3IX count_2181__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i17.GSR = "ENABLED";
    FD1S3IX count_2181__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i18.GSR = "ENABLED";
    FD1S3IX count_2181__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i19.GSR = "ENABLED";
    FD1S3IX count_2181__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i20.GSR = "ENABLED";
    FD1S3IX count_2181__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i21.GSR = "ENABLED";
    FD1S3IX count_2181__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i22.GSR = "ENABLED";
    FD1S3IX count_2181__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i23.GSR = "ENABLED";
    FD1S3IX count_2181__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i24.GSR = "ENABLED";
    FD1S3IX count_2181__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i25.GSR = "ENABLED";
    FD1S3IX count_2181__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i26.GSR = "ENABLED";
    FD1S3IX count_2181__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i27.GSR = "ENABLED";
    FD1S3IX count_2181__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i28.GSR = "ENABLED";
    FD1S3IX count_2181__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i29.GSR = "ENABLED";
    FD1S3IX count_2181__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i30.GSR = "ENABLED";
    FD1S3IX count_2181__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i31.GSR = "ENABLED";
    CCU2D sub_1736_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27535));
    defparam sub_1736_add_2_2.INIT0 = 16'h0000;
    defparam sub_1736_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1736_add_2_2.INJECT1_0 = "NO";
    defparam sub_1736_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27922), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_33.INIT1 = 16'h0000;
    defparam count_2181_add_4_33.INJECT1_0 = "NO";
    defparam count_2181_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27921), .COUT(n27922), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_31.INJECT1_0 = "NO";
    defparam count_2181_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27920), .COUT(n27921), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_29.INJECT1_0 = "NO";
    defparam count_2181_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27919), .COUT(n27920), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_27.INJECT1_0 = "NO";
    defparam count_2181_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27918), .COUT(n27919), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_25.INJECT1_0 = "NO";
    defparam count_2181_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27917), .COUT(n27918), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_23.INJECT1_0 = "NO";
    defparam count_2181_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27916), .COUT(n27917), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_21.INJECT1_0 = "NO";
    defparam count_2181_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27915), .COUT(n27916), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_19.INJECT1_0 = "NO";
    defparam count_2181_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27914), .COUT(n27915), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_17.INJECT1_0 = "NO";
    defparam count_2181_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27913), .COUT(n27914), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_15.INJECT1_0 = "NO";
    defparam count_2181_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27912), .COUT(n27913), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_13.INJECT1_0 = "NO";
    defparam count_2181_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27911), .COUT(n27912), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_11.INJECT1_0 = "NO";
    defparam count_2181_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27910), .COUT(n27911), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_9.INJECT1_0 = "NO";
    defparam count_2181_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27909), .COUT(n27910), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_7.INJECT1_0 = "NO";
    defparam count_2181_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27908), .COUT(n27909), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_5.INJECT1_0 = "NO";
    defparam count_2181_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27907), .COUT(n27908), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_3.INJECT1_0 = "NO";
    defparam count_2181_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27907), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_1.INIT0 = 16'hF000;
    defparam count_2181_add_4_1.INIT1 = 16'h0555;
    defparam count_2181_add_4_1.INJECT1_0 = "NO";
    defparam count_2181_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27550), .S0(n7264));
    defparam sub_1736_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1736_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1736_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1736_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27549), .COUT(n27550));
    defparam sub_1736_add_2_32.INIT0 = 16'h5555;
    defparam sub_1736_add_2_32.INIT1 = 16'h5555;
    defparam sub_1736_add_2_32.INJECT1_0 = "NO";
    defparam sub_1736_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27548), .COUT(n27549));
    defparam sub_1736_add_2_30.INIT0 = 16'h5555;
    defparam sub_1736_add_2_30.INIT1 = 16'h5555;
    defparam sub_1736_add_2_30.INJECT1_0 = "NO";
    defparam sub_1736_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27547), .COUT(n27548));
    defparam sub_1736_add_2_28.INIT0 = 16'h5555;
    defparam sub_1736_add_2_28.INIT1 = 16'h5555;
    defparam sub_1736_add_2_28.INJECT1_0 = "NO";
    defparam sub_1736_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27546), .COUT(n27547));
    defparam sub_1736_add_2_26.INIT0 = 16'h5555;
    defparam sub_1736_add_2_26.INIT1 = 16'h5555;
    defparam sub_1736_add_2_26.INJECT1_0 = "NO";
    defparam sub_1736_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27545), .COUT(n27546));
    defparam sub_1736_add_2_24.INIT0 = 16'h5555;
    defparam sub_1736_add_2_24.INIT1 = 16'h5555;
    defparam sub_1736_add_2_24.INJECT1_0 = "NO";
    defparam sub_1736_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27544), .COUT(n27545));
    defparam sub_1736_add_2_22.INIT0 = 16'h5555;
    defparam sub_1736_add_2_22.INIT1 = 16'h5555;
    defparam sub_1736_add_2_22.INJECT1_0 = "NO";
    defparam sub_1736_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27543), .COUT(n27544));
    defparam sub_1736_add_2_20.INIT0 = 16'h5555;
    defparam sub_1736_add_2_20.INIT1 = 16'h5555;
    defparam sub_1736_add_2_20.INJECT1_0 = "NO";
    defparam sub_1736_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27542), .COUT(n27543));
    defparam sub_1736_add_2_18.INIT0 = 16'h5555;
    defparam sub_1736_add_2_18.INIT1 = 16'h5555;
    defparam sub_1736_add_2_18.INJECT1_0 = "NO";
    defparam sub_1736_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27541), .COUT(n27542));
    defparam sub_1736_add_2_16.INIT0 = 16'h5555;
    defparam sub_1736_add_2_16.INIT1 = 16'h5555;
    defparam sub_1736_add_2_16.INJECT1_0 = "NO";
    defparam sub_1736_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27540), .COUT(n27541));
    defparam sub_1736_add_2_14.INIT0 = 16'h5555;
    defparam sub_1736_add_2_14.INIT1 = 16'h5555;
    defparam sub_1736_add_2_14.INJECT1_0 = "NO";
    defparam sub_1736_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27539), .COUT(n27540));
    defparam sub_1736_add_2_12.INIT0 = 16'h5555;
    defparam sub_1736_add_2_12.INIT1 = 16'h5555;
    defparam sub_1736_add_2_12.INJECT1_0 = "NO";
    defparam sub_1736_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27538), .COUT(n27539));
    defparam sub_1736_add_2_10.INIT0 = 16'h5555;
    defparam sub_1736_add_2_10.INIT1 = 16'h5555;
    defparam sub_1736_add_2_10.INJECT1_0 = "NO";
    defparam sub_1736_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27537), .COUT(n27538));
    defparam sub_1736_add_2_8.INIT0 = 16'h5555;
    defparam sub_1736_add_2_8.INIT1 = 16'h5555;
    defparam sub_1736_add_2_8.INJECT1_0 = "NO";
    defparam sub_1736_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27536), .COUT(n27537));
    defparam sub_1736_add_2_6.INIT0 = 16'h5555;
    defparam sub_1736_add_2_6.INIT1 = 16'h5555;
    defparam sub_1736_add_2_6.INJECT1_0 = "NO";
    defparam sub_1736_add_2_6.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (state, rdata, debug_c_c, n32472, 
            rx_data, n32452, n34346, n29195, \rdata[1] , n183, n32, 
            bclk, debug_c_7, n31583, n32436, n32543, n32542, n32461, 
            n9396_c, n31642, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [5:0]state;
    output [7:0]rdata;
    input debug_c_c;
    input n32472;
    output [7:0]rx_data;
    input n32452;
    input n34346;
    input n29195;
    output \rdata[1] ;
    input n183;
    output n32;
    output bclk;
    output debug_c_7;
    input n31583;
    input n32436;
    input n32543;
    input n32542;
    input n32461;
    input n9396_c;
    input n31642;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n29, n13984, n13985, n21, n17, n29123, n21_adj_7, n23, 
        n28845, n7934, n7936, n29265, baud_reset, n29427, n31576, 
        n7976, n7974, n7972, n7970, n7968, n7966, n7964;
    wire [7:0]rdata_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n7962, n7960, n7958, n7956, n7954, n7952, n7950;
    wire [5:0]n1;
    
    wire n32489, n32544, n4, n31574, n31575, n32491, n4_adj_8, 
        n29183, n11696, n13, n11875, n19, n55, n27990, n56, 
        n2687;
    wire [7:0]n78;
    
    wire n23308, n219, n30509, n30533;
    
    PFUMX i8219 (.BLUT(n29), .ALUT(n13984), .C0(state[0]), .Z(n13985));
    PFUMX i32 (.BLUT(n21), .ALUT(n17), .C0(state[0]), .Z(n29123));
    PFUMX i36 (.BLUT(n21_adj_7), .ALUT(n23), .C0(state[5]), .Z(n28845));
    FD1P3AX rdata_i0_i0 (.D(n7934), .SP(n32472), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n7936), .SP(n32472), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n29265), .CK(debug_c_c), .CD(n32452), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n29427), .CK(debug_c_c), .PD(n32452), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n28845), .CK(debug_c_c), .CD(n32452), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n31576), .CK(debug_c_c), .CD(n32452), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n13985), .CK(debug_c_c), .CD(n34346), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n29123), .CK(debug_c_c), .CD(n34346), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n29195), .CK(debug_c_c), .CD(n34346), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n7976), .SP(n32472), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n7974), .SP(n32472), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n7972), .SP(n32472), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n7970), .SP(n32472), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n7968), .SP(n32472), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n7966), .SP(n32472), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n7964), .SP(n32472), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n7962), .SP(n32472), .CK(debug_c_c), .Q(rdata_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n7960), .SP(n32472), .CK(debug_c_c), .Q(rdata_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n7958), .SP(n32472), .CK(debug_c_c), .Q(rdata_c[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n7956), .SP(n32472), .CK(debug_c_c), .Q(rdata_c[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n7954), .SP(n32472), .CK(debug_c_c), .Q(rdata_c[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n7952), .SP(n32472), .CK(debug_c_c), .Q(rdata_c[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i1 (.D(n7950), .SP(n32472), .CK(debug_c_c), .Q(\rdata[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    LUT4 i21620_4_lut (.A(n183), .B(state[5]), .C(n1[3]), .D(n32), .Z(n29)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21620_4_lut.init = 16'h3111;
    LUT4 i1_4_lut (.A(state[4]), .B(state[3]), .C(state[2]), .D(state[1]), 
         .Z(n32)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heaaa;
    LUT4 i1_2_lut_rep_364 (.A(state[5]), .B(n32), .Z(n32489)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_364.init = 16'h4444;
    LUT4 i1_3_lut_4_lut (.A(state[5]), .B(n32), .C(state[0]), .D(bclk), 
         .Z(n29265)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut.init = 16'hf400;
    LUT4 i1_4_lut_adj_26 (.A(state[5]), .B(state[2]), .C(n183), .D(n32), 
         .Z(n21)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_26.init = 16'h4505;
    LUT4 i1_2_lut_3_lut (.A(state[3]), .B(n32544), .C(state[4]), .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i33_3_lut (.A(state[1]), .B(state[2]), .C(bclk), .Z(n17)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i33_3_lut.init = 16'hc6c6;
    LUT4 n30413_bdd_3_lut_4_lut (.A(state[3]), .B(n32544), .C(bclk), .D(state[4]), 
         .Z(n31574)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n30413_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_8_i4_3_lut_3_lut (.A(state[3]), .B(n32544), .C(bclk), .Z(n1[3])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam mux_8_i4_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i8218_3_lut_3_lut (.A(state[3]), .B(n32544), .C(bclk), .Z(n13984)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i8218_3_lut_3_lut.init = 16'ha6a6;
    PFUMX i24952 (.BLUT(n31575), .ALUT(n31574), .C0(state[0]), .Z(n31576));
    LUT4 i2_4_lut (.A(bclk), .B(n4), .C(state[0]), .D(n32), .Z(n21_adj_7)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'h4840;
    LUT4 i38_4_lut (.A(n183), .B(n32491), .C(state[0]), .D(n4_adj_8), 
         .Z(n23)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i38_4_lut.init = 16'hf535;
    LUT4 i1_2_lut (.A(state[4]), .B(bclk), .Z(n4_adj_8)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut.init = 16'hdddd;
    FD1S3IX drdy_51 (.D(n29183), .CK(debug_c_c), .CD(n34346), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_27 (.A(n11696), .B(rdata[0]), .C(n31583), .D(n13), 
         .Z(n7934)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_27.init = 16'heca0;
    LUT4 i2927_3_lut_rep_419 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n32544)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2927_3_lut_rep_419.init = 16'h8080;
    LUT4 i2_3_lut (.A(state[0]), .B(state[4]), .C(state[5]), .Z(n11696)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i2934_2_lut_rep_366_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n32491)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2934_2_lut_rep_366_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_adj_28 (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_adj_28.init = 16'hefef;
    LUT4 i1_2_lut_adj_29 (.A(state[1]), .B(bclk), .Z(n11875)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_29.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_30 (.A(rdata[0]), .B(rx_data[0]), .C(n32436), .D(n19), 
         .Z(n7936)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_30.init = 16'heca0;
    LUT4 i4_4_lut (.A(n32543), .B(n32542), .C(state[5]), .D(state[0]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    LUT4 i13_4_lut (.A(state[5]), .B(baud_reset), .C(n32461), .D(n9396_c), 
         .Z(n29427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i13_4_lut.init = 16'hceca;
    LUT4 i1_4_lut_4_lut (.A(state[5]), .B(n32461), .C(n9396_c), .D(debug_c_7), 
         .Z(n29183)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_4_lut.init = 16'hfe22;
    LUT4 i1_4_lut_adj_31 (.A(rdata_c[7]), .B(rx_data[7]), .C(n32436), 
         .D(n19), .Z(n7976)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_31.init = 16'heca0;
    LUT4 i1_4_lut_adj_32 (.A(rdata_c[6]), .B(rx_data[6]), .C(n32436), 
         .D(n19), .Z(n7974)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_32.init = 16'heca0;
    LUT4 i1_4_lut_adj_33 (.A(rdata_c[5]), .B(rx_data[5]), .C(n32436), 
         .D(n19), .Z(n7972)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_33.init = 16'heca0;
    LUT4 i1_4_lut_adj_34 (.A(rdata_c[4]), .B(rx_data[4]), .C(n32436), 
         .D(n19), .Z(n7970)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_34.init = 16'heca0;
    LUT4 i1_4_lut_adj_35 (.A(rdata_c[3]), .B(rx_data[3]), .C(n32436), 
         .D(n19), .Z(n7968)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_35.init = 16'heca0;
    LUT4 i1_4_lut_adj_36 (.A(rdata_c[2]), .B(rx_data[2]), .C(n32436), 
         .D(n19), .Z(n7966)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_36.init = 16'heca0;
    LUT4 i1_4_lut_adj_37 (.A(\rdata[1] ), .B(rx_data[1]), .C(n32436), 
         .D(n19), .Z(n7964)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_37.init = 16'heca0;
    LUT4 i1_4_lut_adj_38 (.A(baud_reset), .B(n55), .C(n27990), .D(n56), 
         .Z(n2687)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_38.init = 16'haaba;
    LUT4 n30413_bdd_4_lut (.A(n32489), .B(state[4]), .C(bclk), .D(n32491), 
         .Z(n31575)) /* synthesis lut_function=(!((B (C (D))+!B !(C (D)))+!A)) */ ;
    defparam n30413_bdd_4_lut.init = 16'h2888;
    LUT4 i1_4_lut_adj_39 (.A(n78[7]), .B(rdata_c[7]), .C(n11696), .D(n13), 
         .Z(n7962)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_39.init = 16'heca0;
    LUT4 i3689_4_lut (.A(rdata_c[7]), .B(n9396_c), .C(n23308), .D(n219), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3689_4_lut.init = 16'hcaaa;
    LUT4 i1_2_lut_adj_40 (.A(state[1]), .B(bclk), .Z(n23308)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_40.init = 16'h8888;
    LUT4 i1_2_lut_adj_41 (.A(state[2]), .B(state[3]), .Z(n219)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_41.init = 16'h8888;
    LUT4 i1_4_lut_adj_42 (.A(n78[6]), .B(rdata_c[6]), .C(n11696), .D(n13), 
         .Z(n7960)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_42.init = 16'heca0;
    LUT4 i3691_4_lut (.A(n9396_c), .B(rdata_c[6]), .C(n11875), .D(n219), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3691_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_43 (.A(n78[5]), .B(rdata_c[5]), .C(n11696), .D(n13), 
         .Z(n7958)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_43.init = 16'heca0;
    LUT4 i3693_4_lut (.A(n9396_c), .B(rdata_c[5]), .C(state[1]), .D(n30509), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3693_4_lut.init = 16'hccac;
    LUT4 i1_3_lut (.A(state[2]), .B(state[3]), .C(bclk), .Z(n30509)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut.init = 16'hbfbf;
    LUT4 i1_4_lut_adj_44 (.A(n78[4]), .B(rdata_c[4]), .C(n11696), .D(n13), 
         .Z(n7956)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_44.init = 16'heca0;
    LUT4 i3695_4_lut (.A(n9396_c), .B(rdata_c[4]), .C(state[1]), .D(n30509), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3695_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_45 (.A(n11696), .B(rdata_c[3]), .C(n78[3]), .D(n13), 
         .Z(n7954)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_45.init = 16'heca0;
    LUT4 i3697_4_lut (.A(n9396_c), .B(rdata_c[3]), .C(n23308), .D(n30533), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3697_4_lut.init = 16'hccac;
    LUT4 i1_2_lut_adj_46 (.A(state[3]), .B(state[2]), .Z(n30533)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_adj_46.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_47 (.A(n11696), .B(rdata_c[2]), .C(n78[2]), .D(n13), 
         .Z(n7952)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_47.init = 16'heca0;
    LUT4 i3699_4_lut (.A(n9396_c), .B(rdata_c[2]), .C(n11875), .D(n30533), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3699_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_48 (.A(n11696), .B(\rdata[1] ), .C(n31642), .D(n13), 
         .Z(n7950)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_48.init = 16'heca0;
    \ClockDividerP(factor=12)_U0  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .baud_reset(baud_reset), .n2687(n2687), .n55(n55), .n27990(n27990), 
            .n56(n56), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (bclk, debug_c_c, baud_reset, n2687, 
            n55, n27990, n56, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input baud_reset;
    input n2687;
    output n55;
    output n27990;
    output n56;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7229;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n52, n44, n35, n54, n48, n36, n46, n32, n50, n40, 
        n27566, n27565, n27564, n27563, n27562, n27561, n27560, 
        n27559, n27558, n27557, n27556, n27874, n27555, n27873, 
        n27872, n27554, n27871, n27870, n27553, n27869, n27868, 
        n27552, n27867, n27866, n27551, n27865, n27864, n27863, 
        n27862, n27861, n27860, n27859;
    
    FD1S3IX clk_o_14 (.D(n7229), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2180__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2687), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i0.GSR = "ENABLED";
    FD1S3IX count_2180__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2687), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i1.GSR = "ENABLED";
    FD1S3IX count_2180__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2687), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i2.GSR = "ENABLED";
    FD1S3IX count_2180__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2687), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i3.GSR = "ENABLED";
    FD1S3IX count_2180__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2687), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i4.GSR = "ENABLED";
    FD1S3IX count_2180__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2687), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i5.GSR = "ENABLED";
    FD1S3IX count_2180__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2687), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i6.GSR = "ENABLED";
    FD1S3IX count_2180__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2687), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i7.GSR = "ENABLED";
    FD1S3IX count_2180__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2687), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i8.GSR = "ENABLED";
    FD1S3IX count_2180__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2687), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i9.GSR = "ENABLED";
    FD1S3IX count_2180__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i10.GSR = "ENABLED";
    FD1S3IX count_2180__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i11.GSR = "ENABLED";
    FD1S3IX count_2180__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i12.GSR = "ENABLED";
    FD1S3IX count_2180__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i13.GSR = "ENABLED";
    FD1S3IX count_2180__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i14.GSR = "ENABLED";
    FD1S3IX count_2180__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i15.GSR = "ENABLED";
    FD1S3IX count_2180__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i16.GSR = "ENABLED";
    FD1S3IX count_2180__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i17.GSR = "ENABLED";
    FD1S3IX count_2180__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i18.GSR = "ENABLED";
    FD1S3IX count_2180__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i19.GSR = "ENABLED";
    FD1S3IX count_2180__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i20.GSR = "ENABLED";
    FD1S3IX count_2180__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i21.GSR = "ENABLED";
    FD1S3IX count_2180__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i22.GSR = "ENABLED";
    FD1S3IX count_2180__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i23.GSR = "ENABLED";
    FD1S3IX count_2180__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i24.GSR = "ENABLED";
    FD1S3IX count_2180__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i25.GSR = "ENABLED";
    FD1S3IX count_2180__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i26.GSR = "ENABLED";
    FD1S3IX count_2180__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i27.GSR = "ENABLED";
    FD1S3IX count_2180__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i28.GSR = "ENABLED";
    FD1S3IX count_2180__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i29.GSR = "ENABLED";
    FD1S3IX count_2180__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i30.GSR = "ENABLED";
    FD1S3IX count_2180__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i31.GSR = "ENABLED";
    LUT4 i26_4_lut (.A(count[30]), .B(n52), .C(n44), .D(count[14]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(count[1]), .B(count[3]), .C(count[0]), .Z(n27990)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[12]), .B(n46), .C(n32), .D(count[18]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[24]), .C(count[31]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[16]), .B(count[10]), .C(count[9]), .D(count[17]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[20]), .B(count[5]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[13]), .B(count[22]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[7]), .B(n50), .C(n40), .D(count[11]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[4]), .B(count[6]), .C(count[8]), .D(count[29]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[26]), .B(count[28]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[25]), .B(count[23]), .C(count[2]), .D(count[27]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[19]), .B(count[21]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11_2_lut.init = 16'heeee;
    CCU2D sub_1734_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27566), .S0(n7229));
    defparam sub_1734_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1734_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1734_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1734_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27565), .COUT(n27566));
    defparam sub_1734_add_2_32.INIT0 = 16'h5555;
    defparam sub_1734_add_2_32.INIT1 = 16'h5555;
    defparam sub_1734_add_2_32.INJECT1_0 = "NO";
    defparam sub_1734_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27564), .COUT(n27565));
    defparam sub_1734_add_2_30.INIT0 = 16'h5555;
    defparam sub_1734_add_2_30.INIT1 = 16'h5555;
    defparam sub_1734_add_2_30.INJECT1_0 = "NO";
    defparam sub_1734_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27563), .COUT(n27564));
    defparam sub_1734_add_2_28.INIT0 = 16'h5555;
    defparam sub_1734_add_2_28.INIT1 = 16'h5555;
    defparam sub_1734_add_2_28.INJECT1_0 = "NO";
    defparam sub_1734_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27562), .COUT(n27563));
    defparam sub_1734_add_2_26.INIT0 = 16'h5555;
    defparam sub_1734_add_2_26.INIT1 = 16'h5555;
    defparam sub_1734_add_2_26.INJECT1_0 = "NO";
    defparam sub_1734_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27561), .COUT(n27562));
    defparam sub_1734_add_2_24.INIT0 = 16'h5555;
    defparam sub_1734_add_2_24.INIT1 = 16'h5555;
    defparam sub_1734_add_2_24.INJECT1_0 = "NO";
    defparam sub_1734_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27560), .COUT(n27561));
    defparam sub_1734_add_2_22.INIT0 = 16'h5555;
    defparam sub_1734_add_2_22.INIT1 = 16'h5555;
    defparam sub_1734_add_2_22.INJECT1_0 = "NO";
    defparam sub_1734_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27559), .COUT(n27560));
    defparam sub_1734_add_2_20.INIT0 = 16'h5555;
    defparam sub_1734_add_2_20.INIT1 = 16'h5555;
    defparam sub_1734_add_2_20.INJECT1_0 = "NO";
    defparam sub_1734_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27558), .COUT(n27559));
    defparam sub_1734_add_2_18.INIT0 = 16'h5555;
    defparam sub_1734_add_2_18.INIT1 = 16'h5555;
    defparam sub_1734_add_2_18.INJECT1_0 = "NO";
    defparam sub_1734_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27557), .COUT(n27558));
    defparam sub_1734_add_2_16.INIT0 = 16'h5555;
    defparam sub_1734_add_2_16.INIT1 = 16'h5555;
    defparam sub_1734_add_2_16.INJECT1_0 = "NO";
    defparam sub_1734_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27556), .COUT(n27557));
    defparam sub_1734_add_2_14.INIT0 = 16'h5555;
    defparam sub_1734_add_2_14.INIT1 = 16'h5555;
    defparam sub_1734_add_2_14.INJECT1_0 = "NO";
    defparam sub_1734_add_2_14.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27874), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_33.INIT1 = 16'h0000;
    defparam count_2180_add_4_33.INJECT1_0 = "NO";
    defparam count_2180_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27555), .COUT(n27556));
    defparam sub_1734_add_2_12.INIT0 = 16'h5555;
    defparam sub_1734_add_2_12.INIT1 = 16'h5555;
    defparam sub_1734_add_2_12.INJECT1_0 = "NO";
    defparam sub_1734_add_2_12.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27873), .COUT(n27874), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_31.INJECT1_0 = "NO";
    defparam count_2180_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27872), .COUT(n27873), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_29.INJECT1_0 = "NO";
    defparam count_2180_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27554), .COUT(n27555));
    defparam sub_1734_add_2_10.INIT0 = 16'h5555;
    defparam sub_1734_add_2_10.INIT1 = 16'h5555;
    defparam sub_1734_add_2_10.INJECT1_0 = "NO";
    defparam sub_1734_add_2_10.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27871), .COUT(n27872), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_27.INJECT1_0 = "NO";
    defparam count_2180_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27870), .COUT(n27871), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_25.INJECT1_0 = "NO";
    defparam count_2180_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27553), .COUT(n27554));
    defparam sub_1734_add_2_8.INIT0 = 16'h5555;
    defparam sub_1734_add_2_8.INIT1 = 16'h5555;
    defparam sub_1734_add_2_8.INJECT1_0 = "NO";
    defparam sub_1734_add_2_8.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27869), .COUT(n27870), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_23.INJECT1_0 = "NO";
    defparam count_2180_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27868), .COUT(n27869), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_21.INJECT1_0 = "NO";
    defparam count_2180_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27552), .COUT(n27553));
    defparam sub_1734_add_2_6.INIT0 = 16'h5555;
    defparam sub_1734_add_2_6.INIT1 = 16'h5555;
    defparam sub_1734_add_2_6.INJECT1_0 = "NO";
    defparam sub_1734_add_2_6.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27867), .COUT(n27868), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_19.INJECT1_0 = "NO";
    defparam count_2180_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27866), .COUT(n27867), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_17.INJECT1_0 = "NO";
    defparam count_2180_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27551), .COUT(n27552));
    defparam sub_1734_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1734_add_2_4.INIT1 = 16'h5555;
    defparam sub_1734_add_2_4.INJECT1_0 = "NO";
    defparam sub_1734_add_2_4.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27865), .COUT(n27866), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_15.INJECT1_0 = "NO";
    defparam count_2180_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27864), .COUT(n27865), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_13.INJECT1_0 = "NO";
    defparam count_2180_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27551));
    defparam sub_1734_add_2_2.INIT0 = 16'h0000;
    defparam sub_1734_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1734_add_2_2.INJECT1_0 = "NO";
    defparam sub_1734_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27863), .COUT(n27864), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_11.INJECT1_0 = "NO";
    defparam count_2180_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27862), .COUT(n27863), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_9.INJECT1_0 = "NO";
    defparam count_2180_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27861), .COUT(n27862), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_7.INJECT1_0 = "NO";
    defparam count_2180_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27860), .COUT(n27861), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_5.INJECT1_0 = "NO";
    defparam count_2180_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27859), .COUT(n27860), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_3.INJECT1_0 = "NO";
    defparam count_2180_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27859), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_1.INIT0 = 16'hF000;
    defparam count_2180_add_4_1.INIT1 = 16'h0555;
    defparam count_2180_add_4_1.INJECT1_0 = "NO";
    defparam count_2180_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (GND_net, n224, n32486, n34347, 
            n32387, n32473, n32405, rw, n30450, n32420, n30283, 
            n12434, \register_addr[0] , debug_c_c, n34351, n3451, 
            n34348, \read_size[0] , n11966, n30743, n34349, Stepper_X_M0_c_0, 
            n579, prev_select, n32435, n34350, \register_addr[5] , 
            n34344, n32378, \steps_reg[7] , n30364, limit_c_0, n32509, 
            n32508, n32488, n302, \register_addr[1] , n32527, n32453, 
            read_value, \databus[31] , n34352, \databus[30] , \databus[29] , 
            \databus[26] , \databus[13] , \databus[11] , \databus[10] , 
            \databus[9] , \databus[7] , \databus[6] , \databus[5] , 
            n608, n610, \control_reg[7] , Stepper_X_En_c, n34353, 
            Stepper_X_Dir_c, \databus[3] , Stepper_X_M2_c_2, Stepper_X_M1_c_1, 
            \databus[1] , \read_size[2] , n32463, \register_addr[4] , 
            \register_addr[3] , n11753, n30431, n18, \register_addr[6] , 
            \register_addr[7] , n32478, \databus[8] , \databus[12] , 
            \databus[14] , \databus[15] , \databus[16] , \databus[17] , 
            \databus[18] , \databus[19] , \databus[20] , \databus[21] , 
            \databus[22] , \databus[23] , n32388, n32525, n20291, 
            n28386, \databus[24] , \databus[25] , \databus[27] , \databus[28] , 
            n11645, n32413, n30594, n8048, VCC_net, Stepper_X_nFault_c, 
            Stepper_X_Step_c, n9, n28360) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [31:0]n224;
    input n32486;
    input n34347;
    input n32387;
    input n32473;
    input n32405;
    input rw;
    input n30450;
    input n32420;
    input n30283;
    output n12434;
    input \register_addr[0] ;
    input debug_c_c;
    input n34351;
    input [31:0]n3451;
    input n34348;
    output \read_size[0] ;
    input n11966;
    output n30743;
    input n34349;
    output Stepper_X_M0_c_0;
    input n579;
    output prev_select;
    input n32435;
    input n34350;
    input \register_addr[5] ;
    input n34344;
    output n32378;
    output \steps_reg[7] ;
    input n30364;
    input limit_c_0;
    output n32509;
    input n32508;
    input n32488;
    output n302;
    input \register_addr[1] ;
    input n32527;
    output n32453;
    output [31:0]read_value;
    input \databus[31] ;
    input n34352;
    input \databus[30] ;
    input \databus[29] ;
    input \databus[26] ;
    input \databus[13] ;
    input \databus[11] ;
    input \databus[10] ;
    input \databus[9] ;
    input \databus[7] ;
    input \databus[6] ;
    input \databus[5] ;
    input n608;
    input n610;
    output \control_reg[7] ;
    output Stepper_X_En_c;
    input n34353;
    output Stepper_X_Dir_c;
    input \databus[3] ;
    output Stepper_X_M2_c_2;
    output Stepper_X_M1_c_1;
    input \databus[1] ;
    output \read_size[2] ;
    input n32463;
    input \register_addr[4] ;
    input \register_addr[3] ;
    input n11753;
    output n30431;
    input n18;
    input \register_addr[6] ;
    input \register_addr[7] ;
    output n32478;
    input \databus[8] ;
    input \databus[12] ;
    input \databus[14] ;
    input \databus[15] ;
    input \databus[16] ;
    input \databus[17] ;
    input \databus[18] ;
    input \databus[19] ;
    input \databus[20] ;
    input \databus[21] ;
    input \databus[22] ;
    input \databus[23] ;
    input n32388;
    input n32525;
    input n20291;
    output n28386;
    input \databus[24] ;
    input \databus[25] ;
    input \databus[27] ;
    input \databus[28] ;
    output n11645;
    input n32413;
    output n30594;
    output n8048;
    input VCC_net;
    input Stepper_X_nFault_c;
    output Stepper_X_Step_c;
    input n9;
    output n28360;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27775;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n27776, n12540, n32382, n30895, n30896, n30897, n56, 
        n46, n60, prev_step_clk, step_clk, limit_latched, n182, 
        prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n12480, n30367, n30233, n30371, n30369, n30368, n30366, 
        n30370, n30381, n30380, n30382, n30383, n30384, n30385, 
        n30386, n30387, n30365, n30388, n30372, n32376, n9614;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire fault_latched, n30847, n30848, n1, n2, n1_adj_1, n2_adj_2, 
        n1_adj_3, n2_adj_4, int_step, n11, n32393, n1_adj_5, n2_adj_6, 
        n32495, n27774, n27773, n27772, n27771, n17314, n30856, 
        n30857, n30858, n41, n50, n54, n42, n30849, n52, n38;
    wire [31:0]n5188;
    
    wire n30379, n30378, n30377, n30376, n30375, n30374, n30373, 
        n62, n58, n49, n27786, n27785, n27784, n27783, n27782, 
        n27781, n27780, n27779, n27778, n27777;
    
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27775), .COUT(n27776), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    LUT4 i24744_2_lut_4_lut_4_lut (.A(n32486), .B(n34347), .C(n32387), 
         .D(n32473), .Z(n12540)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i24744_2_lut_4_lut_4_lut.init = 16'hccdc;
    LUT4 i24754_3_lut_rep_257_4_lut_4_lut (.A(n32486), .B(n32473), .C(n32405), 
         .D(rw), .Z(n32382)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i24754_3_lut_rep_257_4_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_4_lut (.A(n30450), .B(n32420), .C(n30283), .D(n34347), 
         .Z(n12434)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff80;
    PFUMX i24539 (.BLUT(n30895), .ALUT(n30896), .C0(\register_addr[0] ), 
          .Z(n30897));
    FD1S3IX steps_reg__i19 (.D(n3451[19]), .CK(debug_c_c), .CD(n34351), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    LUT4 i28_4_lut (.A(steps_reg[2]), .B(n56), .C(n46), .D(steps_reg[16]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    FD1S3IX steps_reg__i18 (.D(n3451[18]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3451[17]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3451[16]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3451[0]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3451[15]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3451[14]), .CK(debug_c_c), .CD(n34348), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n30743), .SP(n11966), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3451[13]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3451[12]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12540), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12480), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3451[11]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32435), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3451[10]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3451[9]), .CK(debug_c_c), .CD(n34349), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3451[8]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_253_3_lut_4_lut (.A(n32435), .B(prev_select), .C(\register_addr[5] ), 
         .D(n34344), .Z(n32378)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_253_3_lut_4_lut.init = 16'h0002;
    FD1S3IX steps_reg__i7 (.D(n3451[7]), .CK(debug_c_c), .CD(n34350), 
            .Q(\steps_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3451[6]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(div_factor_reg[18]), .B(n30364), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n30367)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 equal_138_i16_1_lut_2_lut_3_lut_4_lut (.A(n32509), .B(n32508), 
         .C(n32488), .D(\register_addr[0] ), .Z(n302)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_138_i16_1_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32509), .B(n32508), .C(\register_addr[1] ), 
         .D(n32527), .Z(n30233)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1S3IX steps_reg__i5 (.D(n3451[5]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3451[4]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3451[3]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    LUT4 i24833_2_lut_3_lut_4_lut (.A(n32509), .B(n32508), .C(\register_addr[1] ), 
         .D(n32527), .Z(n30743)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i24833_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 equal_138_i15_2_lut_rep_328_3_lut_4_lut (.A(n32509), .B(n32508), 
         .C(n32488), .D(\register_addr[0] ), .Z(n32453)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_138_i15_2_lut_rep_328_3_lut_4_lut.init = 16'hfffe;
    FD1S3IX steps_reg__i2 (.D(n3451[2]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3451[1]), .CK(debug_c_c), .CD(n34350), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n30371), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n30369), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n30367), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30368), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30366), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30370), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30381), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30380), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30382), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n30383), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n30384), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30385), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30386), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30387), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30365), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n30388), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_1 (.A(div_factor_reg[15]), .B(n30364), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n30372)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_1.init = 16'hc088;
    FD1P3IX div_factor_reg_i31 (.D(\databus[31] ), .SP(n32376), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(\databus[30] ), .SP(n32376), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(\databus[29] ), .SP(n32376), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(\databus[26] ), .SP(n32376), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(\databus[13] ), .SP(n32376), .PD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(\databus[11] ), .SP(n32376), .PD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(\databus[10] ), .SP(n32376), .PD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(\databus[9] ), .SP(n32376), .PD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(\databus[7] ), .SP(n32376), .PD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(\databus[6] ), .SP(n32376), .PD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(\databus[5] ), .SP(n32376), .PD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n12480), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12480), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(\databus[7] ), .SP(n32382), .CD(n9614), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(\databus[6] ), .SP(n32382), .PD(n34353), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(\databus[5] ), .SP(n32382), .PD(n34353), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n12540), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(\databus[3] ), .SP(n32382), .PD(n34353), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n12540), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(\databus[1] ), .SP(n32382), .PD(n34353), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n30233), .SP(n11966), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3451[31]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3451[30]), .CK(debug_c_c), .CD(n34353), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3451[29]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3451[28]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3451[27]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3451[26]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3451[25]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3451[24]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3451[23]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3451[22]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3451[21]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3451[20]), .CK(debug_c_c), .CD(n32463), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    LUT4 i24489_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30847)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24489_3_lut.init = 16'hcaca;
    LUT4 i24490_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24490_3_lut.init = 16'hcaca;
    LUT4 i14226_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14226_2_lut.init = 16'h2222;
    LUT4 mux_1600_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1600_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i14225_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14225_2_lut.init = 16'h2222;
    LUT4 mux_1600_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2_adj_2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1600_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 i14224_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_3)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14224_2_lut.init = 16'h2222;
    LUT4 mux_1600_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2_adj_4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1600_Mux_5_i2_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n32393), .SP(n11), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i14223_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_5)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14223_2_lut.init = 16'h2222;
    LUT4 mux_1600_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1600_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 i14240_2_lut_rep_370 (.A(\register_addr[4] ), .B(\register_addr[3] ), 
         .Z(n32495)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14240_2_lut_rep_370.init = 16'heeee;
    LUT4 i1_4_lut_adj_2 (.A(div_factor_reg[24]), .B(n30364), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n30382)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_2.init = 16'hc088;
    LUT4 i1_4_lut_adj_3 (.A(div_factor_reg[25]), .B(n30364), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n30383)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_3.init = 16'hc088;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[4] ), .B(\register_addr[3] ), 
         .C(n11753), .Z(n30431)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_4_lut_adj_4 (.A(div_factor_reg[26]), .B(n30364), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n30384)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_4.init = 16'hc088;
    CCU2D sub_125_add_2_9 (.A0(\steps_reg[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27774), .COUT(n27775), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27773), .COUT(n27774), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27772), .COUT(n27773), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_5 (.A(div_factor_reg[27]), .B(n30364), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n30385)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_5.init = 16'hc088;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27771), .COUT(n27772), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n18), .D1(prev_step_clk), 
          .COUT(n27771), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_6 (.A(div_factor_reg[28]), .B(n30364), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n30386)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_6.init = 16'hc088;
    LUT4 i1_4_lut_adj_7 (.A(div_factor_reg[29]), .B(n30364), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n30387)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_7.init = 16'hc088;
    LUT4 i1_4_lut_adj_8 (.A(div_factor_reg[30]), .B(n30364), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n30365)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_8.init = 16'hc088;
    LUT4 i1_4_lut_adj_9 (.A(div_factor_reg[31]), .B(n30364), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n30388)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_9.init = 16'hc088;
    LUT4 i1_4_lut_adj_10 (.A(div_factor_reg[19]), .B(n30364), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n30368)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_10.init = 16'hc088;
    LUT4 i11563_3_lut (.A(\control_reg[7] ), .B(div_factor_reg[7]), .C(\register_addr[1] ), 
         .Z(n17314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11563_3_lut.init = 16'hcaca;
    LUT4 i3853_3_lut (.A(prev_limit_latched), .B(n34347), .C(limit_latched), 
         .Z(n9614)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3853_3_lut.init = 16'hdcdc;
    LUT4 equal_138_i13_2_lut_rep_384 (.A(\register_addr[6] ), .B(\register_addr[7] ), 
         .Z(n32509)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_138_i13_2_lut_rep_384.init = 16'heeee;
    LUT4 i1_2_lut_rep_353_3_lut_4_lut (.A(\register_addr[6] ), .B(\register_addr[7] ), 
         .C(\register_addr[5] ), .D(\register_addr[4] ), .Z(n32478)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_353_3_lut_4_lut.init = 16'hfffe;
    PFUMX i24500 (.BLUT(n30856), .ALUT(n30857), .C0(\register_addr[1] ), 
          .Z(n30858));
    FD1P3IX div_factor_reg_i1 (.D(\databus[1] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(\databus[3] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(\steps_reg[7] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(steps_reg[20]), .B(steps_reg[21]), .C(steps_reg[11]), 
         .D(steps_reg[25]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[6]), .C(steps_reg[5]), 
         .D(steps_reg[10]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_11 (.A(div_factor_reg[20]), .B(n30364), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n30366)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_11.init = 16'hc088;
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    FD1P3IX div_factor_reg_i8 (.D(\databus[8] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(\databus[12] ), .SP(n12480), .CD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(\databus[14] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_12 (.A(div_factor_reg[21]), .B(n30364), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n30370)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_12.init = 16'hc088;
    LUT4 i1_4_lut_adj_13 (.A(div_factor_reg[22]), .B(n30364), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n30381)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_13.init = 16'hc088;
    FD1P3IX div_factor_reg_i15 (.D(\databus[15] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    LUT4 i24_4_lut (.A(steps_reg[29]), .B(steps_reg[3]), .C(steps_reg[13]), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    FD1P3IX div_factor_reg_i16 (.D(\databus[16] ), .SP(n12480), .CD(n34351), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_14 (.A(div_factor_reg[23]), .B(n30364), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n30380)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_14.init = 16'hc088;
    FD1P3IX div_factor_reg_i17 (.D(\databus[17] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(\databus[18] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(\databus[19] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(\databus[20] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(\databus[21] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(\databus[22] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    LUT4 i14_2_lut (.A(steps_reg[15]), .B(steps_reg[23]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    FD1P3IX div_factor_reg_i23 (.D(\databus[23] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30849), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i20_4_lut (.A(steps_reg[1]), .B(steps_reg[4]), .C(steps_reg[0]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    FD1P3IX read_value__i2 (.D(n30897), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    LUT4 i24782_4_lut (.A(n32525), .B(n20291), .C(\register_addr[5] ), 
         .D(n32495), .Z(n28386)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24782_4_lut.init = 16'h0001;
    LUT4 i6_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    FD1P3IX read_value__i3 (.D(n5188[3]), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(\databus[24] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5188[4]), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(\databus[25] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n5188[5]), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(\databus[27] ), .SP(n12480), .CD(n34348), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n5188[6]), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(\databus[28] ), .SP(n12480), .CD(n34352), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n5188[7]), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30379), .SP(n11966), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n30378), .SP(n11966), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n30377), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n11645)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i2_4_lut (.A(n32478), .B(n32413), .C(n32527), .D(n30594), .Z(n8048)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0400;
    LUT4 i24241_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n30594)) /* synthesis lut_function=(A (B)) */ ;
    defparam i24241_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_15 (.A(n30450), .B(\register_addr[4] ), .C(n32378), 
         .D(n34347), .Z(n12480)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_15.init = 16'hff20;
    FD1P3AX read_value__i11 (.D(n30376), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30375), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30374), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30373), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_251_4_lut (.A(\register_addr[5] ), .B(n32387), .C(\register_addr[4] ), 
         .D(n30450), .Z(n32376)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_rep_251_4_lut.init = 16'h0400;
    FD1P3IX read_value__i0 (.D(n30858), .SP(n11966), .CD(n32388), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n30372), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[26]), .B(n52), .C(n38), .D(steps_reg[9]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i24498_3_lut (.A(Stepper_X_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24498_3_lut.init = 16'hcaca;
    LUT4 i24499_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24499_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_16 (.A(div_factor_reg[8]), .B(n30364), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n30379)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_16.init = 16'hc088;
    PFUMX i24491 (.BLUT(n30847), .ALUT(n30848), .C0(\register_addr[1] ), 
          .Z(n30849));
    LUT4 i1_2_lut_adj_17 (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_17.init = 16'h9999;
    LUT4 i1_4_lut_adj_18 (.A(div_factor_reg[9]), .B(n30364), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n30378)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_18.init = 16'hc088;
    LUT4 i24537_3_lut (.A(Stepper_X_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24537_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_19 (.A(div_factor_reg[10]), .B(n30364), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n30377)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_19.init = 16'hc088;
    PFUMX mux_1600_Mux_3_i3 (.BLUT(n1), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n5188[3]));
    PFUMX mux_1600_Mux_4_i3 (.BLUT(n1_adj_1), .ALUT(n2_adj_2), .C0(\register_addr[1] ), 
          .Z(n5188[4]));
    LUT4 i24538_3_lut (.A(n18), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24538_3_lut.init = 16'hcaca;
    PFUMX mux_1600_Mux_5_i3 (.BLUT(n1_adj_3), .ALUT(n2_adj_4), .C0(\register_addr[1] ), 
          .Z(n5188[5]));
    PFUMX mux_1600_Mux_6_i3 (.BLUT(n1_adj_5), .ALUT(n2_adj_6), .C0(\register_addr[1] ), 
          .Z(n5188[6]));
    PFUMX i11565 (.BLUT(n17314), .ALUT(n9), .C0(\register_addr[0] ), .Z(n5188[7]));
    LUT4 i1_4_lut_adj_20 (.A(div_factor_reg[11]), .B(n30364), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n30376)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_20.init = 16'hc088;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28360)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_21 (.A(div_factor_reg[12]), .B(n30364), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n30375)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_21.init = 16'hc088;
    LUT4 i1_4_lut_adj_22 (.A(div_factor_reg[13]), .B(n30364), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n30374)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_22.init = 16'hc088;
    LUT4 i17_4_lut (.A(steps_reg[24]), .B(steps_reg[18]), .C(steps_reg[28]), 
         .D(steps_reg[8]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_23 (.A(div_factor_reg[14]), .B(n30364), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n30373)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_23.init = 16'hc088;
    LUT4 i1_4_lut_adj_24 (.A(div_factor_reg[16]), .B(n30364), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n30371)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_24.init = 16'hc088;
    LUT4 i1_4_lut_adj_25 (.A(div_factor_reg[17]), .B(n30364), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n30369)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_25.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27786), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27785), .COUT(n27786), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27784), .COUT(n27785), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27783), .COUT(n27784), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27782), .COUT(n27783), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27781), .COUT(n27782), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27780), .COUT(n27781), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27779), .COUT(n27780), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27778), .COUT(n27779), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27777), .COUT(n27778), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27776), .COUT(n27777), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    ClockDivider_U8 step_clk_gen (.n34347(n34347), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n32463(n32463), .prev_step_clk(prev_step_clk), 
            .n18(n18), .n32393(n32393), .n11(n11), .GND_net(GND_net), 
            .div_factor_reg({div_factor_reg})) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (n34347, step_clk, debug_c_c, n32463, prev_step_clk, 
            n18, n32393, n11, GND_net, div_factor_reg) /* synthesis syn_module_defined=1 */ ;
    input n34347;
    output step_clk;
    input debug_c_c;
    input n32463;
    input prev_step_clk;
    input n18;
    output n32393;
    output n11;
    input GND_net;
    input [31:0]div_factor_reg;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n6848, n32370, n6882, n14150, n6813;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27722;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n27721, n27720, n27719, n27718, n27717, n27716, n27715, 
        n27714, n27713, n27712, n27711, n27710, n27709, n27708, 
        n27707, n27534, n27533, n27532, n27531, n27530, n27529, 
        n27528, n27527, n27526, n27525, n27524, n27523, n27522, 
        n27521, n27520, n27519, n27518, n27517, n27516, n27515, 
        n27514, n27513, n27512, n27511, n27510, n27509, n27508, 
        n27507, n27506, n27505, n27504, n27503, n27502, n27501, 
        n27500, n27499, n27498, n27497, n27496, n27495, n27494, 
        n27493, n27492, n27491, n27490, n27489, n27488, n27487, 
        n27890, n27889, n27888, n27887, n27886, n27885, n27884, 
        n27883, n27882, n27881, n27880, n27879, n27878, n27877, 
        n27876, n27875;
    
    LUT4 i954_2_lut_rep_245 (.A(n6848), .B(n34347), .Z(n32370)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i954_2_lut_rep_245.init = 16'heeee;
    LUT4 i8470_2_lut_3_lut (.A(n6848), .B(n34347), .C(n6882), .Z(n14150)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8470_2_lut_3_lut.init = 16'he0e0;
    FD1S3IX clk_o_22 (.D(n6813), .CK(debug_c_c), .CD(n32463), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2176__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i0.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_268 (.A(prev_step_clk), .B(n18), .C(step_clk), .Z(n32393)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i2_3_lut_rep_268.init = 16'h4040;
    LUT4 i1_4_lut_4_lut (.A(prev_step_clk), .B(n18), .C(step_clk), .D(n34347), 
         .Z(n11)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i1_4_lut_4_lut.init = 16'h004a;
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27722), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27721), .COUT(n27722), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27720), .COUT(n27721), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27719), .COUT(n27720), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27718), .COUT(n27719), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27717), .COUT(n27718), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27716), .COUT(n27717), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27715), .COUT(n27716), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27714), .COUT(n27715), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27713), .COUT(n27714), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32370), .PD(n14150), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27712), .COUT(n27713), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27711), .COUT(n27712), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    FD1S3IX count_2176__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27710), .COUT(n27711), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    FD1S3IX count_2176__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i2.GSR = "ENABLED";
    FD1S3IX count_2176__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i3.GSR = "ENABLED";
    FD1S3IX count_2176__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i4.GSR = "ENABLED";
    FD1S3IX count_2176__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i5.GSR = "ENABLED";
    FD1S3IX count_2176__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i6.GSR = "ENABLED";
    FD1S3IX count_2176__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i7.GSR = "ENABLED";
    FD1S3IX count_2176__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i8.GSR = "ENABLED";
    FD1S3IX count_2176__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i9.GSR = "ENABLED";
    FD1S3IX count_2176__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i10.GSR = "ENABLED";
    FD1S3IX count_2176__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i11.GSR = "ENABLED";
    FD1S3IX count_2176__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i12.GSR = "ENABLED";
    FD1S3IX count_2176__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i13.GSR = "ENABLED";
    FD1S3IX count_2176__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i14.GSR = "ENABLED";
    FD1S3IX count_2176__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i15.GSR = "ENABLED";
    FD1S3IX count_2176__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i16.GSR = "ENABLED";
    FD1S3IX count_2176__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i17.GSR = "ENABLED";
    FD1S3IX count_2176__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i18.GSR = "ENABLED";
    FD1S3IX count_2176__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i19.GSR = "ENABLED";
    FD1S3IX count_2176__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i20.GSR = "ENABLED";
    FD1S3IX count_2176__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i21.GSR = "ENABLED";
    FD1S3IX count_2176__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i22.GSR = "ENABLED";
    FD1S3IX count_2176__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i23.GSR = "ENABLED";
    FD1S3IX count_2176__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i24.GSR = "ENABLED";
    FD1S3IX count_2176__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i25.GSR = "ENABLED";
    FD1S3IX count_2176__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i26.GSR = "ENABLED";
    FD1S3IX count_2176__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i27.GSR = "ENABLED";
    FD1S3IX count_2176__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i28.GSR = "ENABLED";
    FD1S3IX count_2176__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i29.GSR = "ENABLED";
    FD1S3IX count_2176__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i30.GSR = "ENABLED";
    FD1S3IX count_2176__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32370), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27709), .COUT(n27710), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27708), .COUT(n27709), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27707), .COUT(n27708), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27534), .S1(n6813));
    defparam sub_1714_add_2_33.INIT0 = 16'h5555;
    defparam sub_1714_add_2_33.INIT1 = 16'h0000;
    defparam sub_1714_add_2_33.INJECT1_0 = "NO";
    defparam sub_1714_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27533), .COUT(n27534));
    defparam sub_1714_add_2_31.INIT0 = 16'h5999;
    defparam sub_1714_add_2_31.INIT1 = 16'h5999;
    defparam sub_1714_add_2_31.INJECT1_0 = "NO";
    defparam sub_1714_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27707), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27532), .COUT(n27533));
    defparam sub_1714_add_2_29.INIT0 = 16'h5999;
    defparam sub_1714_add_2_29.INIT1 = 16'h5999;
    defparam sub_1714_add_2_29.INJECT1_0 = "NO";
    defparam sub_1714_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27531), .COUT(n27532));
    defparam sub_1714_add_2_27.INIT0 = 16'h5999;
    defparam sub_1714_add_2_27.INIT1 = 16'h5999;
    defparam sub_1714_add_2_27.INJECT1_0 = "NO";
    defparam sub_1714_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27530), .COUT(n27531));
    defparam sub_1714_add_2_25.INIT0 = 16'h5999;
    defparam sub_1714_add_2_25.INIT1 = 16'h5999;
    defparam sub_1714_add_2_25.INJECT1_0 = "NO";
    defparam sub_1714_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27529), .COUT(n27530));
    defparam sub_1714_add_2_23.INIT0 = 16'h5999;
    defparam sub_1714_add_2_23.INIT1 = 16'h5999;
    defparam sub_1714_add_2_23.INJECT1_0 = "NO";
    defparam sub_1714_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27528), .COUT(n27529));
    defparam sub_1714_add_2_21.INIT0 = 16'h5999;
    defparam sub_1714_add_2_21.INIT1 = 16'h5999;
    defparam sub_1714_add_2_21.INJECT1_0 = "NO";
    defparam sub_1714_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27527), .COUT(n27528));
    defparam sub_1714_add_2_19.INIT0 = 16'h5999;
    defparam sub_1714_add_2_19.INIT1 = 16'h5999;
    defparam sub_1714_add_2_19.INJECT1_0 = "NO";
    defparam sub_1714_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27526), .COUT(n27527));
    defparam sub_1714_add_2_17.INIT0 = 16'h5999;
    defparam sub_1714_add_2_17.INIT1 = 16'h5999;
    defparam sub_1714_add_2_17.INJECT1_0 = "NO";
    defparam sub_1714_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27525), .COUT(n27526));
    defparam sub_1714_add_2_15.INIT0 = 16'h5999;
    defparam sub_1714_add_2_15.INIT1 = 16'h5999;
    defparam sub_1714_add_2_15.INJECT1_0 = "NO";
    defparam sub_1714_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27524), .COUT(n27525));
    defparam sub_1714_add_2_13.INIT0 = 16'h5999;
    defparam sub_1714_add_2_13.INIT1 = 16'h5999;
    defparam sub_1714_add_2_13.INJECT1_0 = "NO";
    defparam sub_1714_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27523), .COUT(n27524));
    defparam sub_1714_add_2_11.INIT0 = 16'h5999;
    defparam sub_1714_add_2_11.INIT1 = 16'h5999;
    defparam sub_1714_add_2_11.INJECT1_0 = "NO";
    defparam sub_1714_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27522), .COUT(n27523));
    defparam sub_1714_add_2_9.INIT0 = 16'h5999;
    defparam sub_1714_add_2_9.INIT1 = 16'h5999;
    defparam sub_1714_add_2_9.INJECT1_0 = "NO";
    defparam sub_1714_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27521), .COUT(n27522));
    defparam sub_1714_add_2_7.INIT0 = 16'h5999;
    defparam sub_1714_add_2_7.INIT1 = 16'h5999;
    defparam sub_1714_add_2_7.INJECT1_0 = "NO";
    defparam sub_1714_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27520), .COUT(n27521));
    defparam sub_1714_add_2_5.INIT0 = 16'h5999;
    defparam sub_1714_add_2_5.INIT1 = 16'h5999;
    defparam sub_1714_add_2_5.INJECT1_0 = "NO";
    defparam sub_1714_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27519), .COUT(n27520));
    defparam sub_1714_add_2_3.INIT0 = 16'h5999;
    defparam sub_1714_add_2_3.INIT1 = 16'h5999;
    defparam sub_1714_add_2_3.INJECT1_0 = "NO";
    defparam sub_1714_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27519));
    defparam sub_1714_add_2_1.INIT0 = 16'h0000;
    defparam sub_1714_add_2_1.INIT1 = 16'h5999;
    defparam sub_1714_add_2_1.INJECT1_0 = "NO";
    defparam sub_1714_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27518), .S1(n6848));
    defparam sub_1716_add_2_33.INIT0 = 16'h5999;
    defparam sub_1716_add_2_33.INIT1 = 16'h0000;
    defparam sub_1716_add_2_33.INJECT1_0 = "NO";
    defparam sub_1716_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27517), .COUT(n27518));
    defparam sub_1716_add_2_31.INIT0 = 16'h5999;
    defparam sub_1716_add_2_31.INIT1 = 16'h5999;
    defparam sub_1716_add_2_31.INJECT1_0 = "NO";
    defparam sub_1716_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    CCU2D sub_1716_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27516), .COUT(n27517));
    defparam sub_1716_add_2_29.INIT0 = 16'h5999;
    defparam sub_1716_add_2_29.INIT1 = 16'h5999;
    defparam sub_1716_add_2_29.INJECT1_0 = "NO";
    defparam sub_1716_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27515), .COUT(n27516));
    defparam sub_1716_add_2_27.INIT0 = 16'h5999;
    defparam sub_1716_add_2_27.INIT1 = 16'h5999;
    defparam sub_1716_add_2_27.INJECT1_0 = "NO";
    defparam sub_1716_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27514), .COUT(n27515));
    defparam sub_1716_add_2_25.INIT0 = 16'h5999;
    defparam sub_1716_add_2_25.INIT1 = 16'h5999;
    defparam sub_1716_add_2_25.INJECT1_0 = "NO";
    defparam sub_1716_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27513), .COUT(n27514));
    defparam sub_1716_add_2_23.INIT0 = 16'h5999;
    defparam sub_1716_add_2_23.INIT1 = 16'h5999;
    defparam sub_1716_add_2_23.INJECT1_0 = "NO";
    defparam sub_1716_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27512), .COUT(n27513));
    defparam sub_1716_add_2_21.INIT0 = 16'h5999;
    defparam sub_1716_add_2_21.INIT1 = 16'h5999;
    defparam sub_1716_add_2_21.INJECT1_0 = "NO";
    defparam sub_1716_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27511), .COUT(n27512));
    defparam sub_1716_add_2_19.INIT0 = 16'h5999;
    defparam sub_1716_add_2_19.INIT1 = 16'h5999;
    defparam sub_1716_add_2_19.INJECT1_0 = "NO";
    defparam sub_1716_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27510), .COUT(n27511));
    defparam sub_1716_add_2_17.INIT0 = 16'h5999;
    defparam sub_1716_add_2_17.INIT1 = 16'h5999;
    defparam sub_1716_add_2_17.INJECT1_0 = "NO";
    defparam sub_1716_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27509), .COUT(n27510));
    defparam sub_1716_add_2_15.INIT0 = 16'h5999;
    defparam sub_1716_add_2_15.INIT1 = 16'h5999;
    defparam sub_1716_add_2_15.INJECT1_0 = "NO";
    defparam sub_1716_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27508), .COUT(n27509));
    defparam sub_1716_add_2_13.INIT0 = 16'h5999;
    defparam sub_1716_add_2_13.INIT1 = 16'h5999;
    defparam sub_1716_add_2_13.INJECT1_0 = "NO";
    defparam sub_1716_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27507), .COUT(n27508));
    defparam sub_1716_add_2_11.INIT0 = 16'h5999;
    defparam sub_1716_add_2_11.INIT1 = 16'h5999;
    defparam sub_1716_add_2_11.INJECT1_0 = "NO";
    defparam sub_1716_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27506), .COUT(n27507));
    defparam sub_1716_add_2_9.INIT0 = 16'h5999;
    defparam sub_1716_add_2_9.INIT1 = 16'h5999;
    defparam sub_1716_add_2_9.INJECT1_0 = "NO";
    defparam sub_1716_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27505), .COUT(n27506));
    defparam sub_1716_add_2_7.INIT0 = 16'h5999;
    defparam sub_1716_add_2_7.INIT1 = 16'h5999;
    defparam sub_1716_add_2_7.INJECT1_0 = "NO";
    defparam sub_1716_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27504), .COUT(n27505));
    defparam sub_1716_add_2_5.INIT0 = 16'h5999;
    defparam sub_1716_add_2_5.INIT1 = 16'h5999;
    defparam sub_1716_add_2_5.INJECT1_0 = "NO";
    defparam sub_1716_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27503), .COUT(n27504));
    defparam sub_1716_add_2_3.INIT0 = 16'h5999;
    defparam sub_1716_add_2_3.INIT1 = 16'h5999;
    defparam sub_1716_add_2_3.INJECT1_0 = "NO";
    defparam sub_1716_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    CCU2D sub_1716_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27503));
    defparam sub_1716_add_2_1.INIT0 = 16'h0000;
    defparam sub_1716_add_2_1.INIT1 = 16'h5999;
    defparam sub_1716_add_2_1.INJECT1_0 = "NO";
    defparam sub_1716_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27502), .S1(n6882));
    defparam sub_1717_add_2_33.INIT0 = 16'hf555;
    defparam sub_1717_add_2_33.INIT1 = 16'h0000;
    defparam sub_1717_add_2_33.INJECT1_0 = "NO";
    defparam sub_1717_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27501), .COUT(n27502));
    defparam sub_1717_add_2_31.INIT0 = 16'hf555;
    defparam sub_1717_add_2_31.INIT1 = 16'hf555;
    defparam sub_1717_add_2_31.INJECT1_0 = "NO";
    defparam sub_1717_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27500), .COUT(n27501));
    defparam sub_1717_add_2_29.INIT0 = 16'hf555;
    defparam sub_1717_add_2_29.INIT1 = 16'hf555;
    defparam sub_1717_add_2_29.INJECT1_0 = "NO";
    defparam sub_1717_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27499), .COUT(n27500));
    defparam sub_1717_add_2_27.INIT0 = 16'hf555;
    defparam sub_1717_add_2_27.INIT1 = 16'hf555;
    defparam sub_1717_add_2_27.INJECT1_0 = "NO";
    defparam sub_1717_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27498), .COUT(n27499));
    defparam sub_1717_add_2_25.INIT0 = 16'hf555;
    defparam sub_1717_add_2_25.INIT1 = 16'hf555;
    defparam sub_1717_add_2_25.INJECT1_0 = "NO";
    defparam sub_1717_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27497), .COUT(n27498));
    defparam sub_1717_add_2_23.INIT0 = 16'hf555;
    defparam sub_1717_add_2_23.INIT1 = 16'hf555;
    defparam sub_1717_add_2_23.INJECT1_0 = "NO";
    defparam sub_1717_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27496), .COUT(n27497));
    defparam sub_1717_add_2_21.INIT0 = 16'hf555;
    defparam sub_1717_add_2_21.INIT1 = 16'hf555;
    defparam sub_1717_add_2_21.INJECT1_0 = "NO";
    defparam sub_1717_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27495), .COUT(n27496));
    defparam sub_1717_add_2_19.INIT0 = 16'hf555;
    defparam sub_1717_add_2_19.INIT1 = 16'hf555;
    defparam sub_1717_add_2_19.INJECT1_0 = "NO";
    defparam sub_1717_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27494), .COUT(n27495));
    defparam sub_1717_add_2_17.INIT0 = 16'hf555;
    defparam sub_1717_add_2_17.INIT1 = 16'hf555;
    defparam sub_1717_add_2_17.INJECT1_0 = "NO";
    defparam sub_1717_add_2_17.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    CCU2D sub_1717_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27493), .COUT(n27494));
    defparam sub_1717_add_2_15.INIT0 = 16'hf555;
    defparam sub_1717_add_2_15.INIT1 = 16'hf555;
    defparam sub_1717_add_2_15.INJECT1_0 = "NO";
    defparam sub_1717_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27492), .COUT(n27493));
    defparam sub_1717_add_2_13.INIT0 = 16'hf555;
    defparam sub_1717_add_2_13.INIT1 = 16'hf555;
    defparam sub_1717_add_2_13.INJECT1_0 = "NO";
    defparam sub_1717_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27491), .COUT(n27492));
    defparam sub_1717_add_2_11.INIT0 = 16'hf555;
    defparam sub_1717_add_2_11.INIT1 = 16'hf555;
    defparam sub_1717_add_2_11.INJECT1_0 = "NO";
    defparam sub_1717_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27490), .COUT(n27491));
    defparam sub_1717_add_2_9.INIT0 = 16'hf555;
    defparam sub_1717_add_2_9.INIT1 = 16'hf555;
    defparam sub_1717_add_2_9.INJECT1_0 = "NO";
    defparam sub_1717_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27489), .COUT(n27490));
    defparam sub_1717_add_2_7.INIT0 = 16'hf555;
    defparam sub_1717_add_2_7.INIT1 = 16'hf555;
    defparam sub_1717_add_2_7.INJECT1_0 = "NO";
    defparam sub_1717_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27488), .COUT(n27489));
    defparam sub_1717_add_2_5.INIT0 = 16'hf555;
    defparam sub_1717_add_2_5.INIT1 = 16'hf555;
    defparam sub_1717_add_2_5.INJECT1_0 = "NO";
    defparam sub_1717_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27487), .COUT(n27488));
    defparam sub_1717_add_2_3.INIT0 = 16'hf555;
    defparam sub_1717_add_2_3.INIT1 = 16'hf555;
    defparam sub_1717_add_2_3.INJECT1_0 = "NO";
    defparam sub_1717_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27487));
    defparam sub_1717_add_2_1.INIT0 = 16'h0000;
    defparam sub_1717_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1717_add_2_1.INJECT1_0 = "NO";
    defparam sub_1717_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32370), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    CCU2D count_2176_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27890), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_33.INIT1 = 16'h0000;
    defparam count_2176_add_4_33.INJECT1_0 = "NO";
    defparam count_2176_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27889), .COUT(n27890), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_31.INJECT1_0 = "NO";
    defparam count_2176_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27888), .COUT(n27889), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_29.INJECT1_0 = "NO";
    defparam count_2176_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27887), .COUT(n27888), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_27.INJECT1_0 = "NO";
    defparam count_2176_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27886), .COUT(n27887), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_25.INJECT1_0 = "NO";
    defparam count_2176_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27885), .COUT(n27886), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_23.INJECT1_0 = "NO";
    defparam count_2176_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27884), .COUT(n27885), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_21.INJECT1_0 = "NO";
    defparam count_2176_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27883), .COUT(n27884), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_19.INJECT1_0 = "NO";
    defparam count_2176_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27882), .COUT(n27883), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_17.INJECT1_0 = "NO";
    defparam count_2176_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27881), .COUT(n27882), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_15.INJECT1_0 = "NO";
    defparam count_2176_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27880), .COUT(n27881), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_13.INJECT1_0 = "NO";
    defparam count_2176_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27879), .COUT(n27880), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_11.INJECT1_0 = "NO";
    defparam count_2176_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27878), .COUT(n27879), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_9.INJECT1_0 = "NO";
    defparam count_2176_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27877), .COUT(n27878), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_7.INJECT1_0 = "NO";
    defparam count_2176_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27876), .COUT(n27877), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_5.INJECT1_0 = "NO";
    defparam count_2176_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27875), .COUT(n27876), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_3.INJECT1_0 = "NO";
    defparam count_2176_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27875), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_1.INIT0 = 16'hF000;
    defparam count_2176_add_4_1.INIT1 = 16'h0555;
    defparam count_2176_add_4_1.INJECT1_0 = "NO";
    defparam count_2176_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (debug_c_c, n241, n34347, n6674, n32375, n31079, 
            n32374, n30942, n12030, n31025, n12031, n30958, n28331, 
            n30940, n28339, n31033, n28345, n31041, n28337, n31057, 
            n28352, n988, n6, n30999, n12138, n31050, n11987, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n241;
    input n34347;
    output n6674;
    output n32375;
    input n31079;
    output n32374;
    input n30942;
    output n12030;
    input n31025;
    output n12031;
    input n30958;
    output n28331;
    input n30940;
    output n28339;
    input n31033;
    output n28345;
    input n31041;
    output n28337;
    input n31057;
    output n28352;
    input n988;
    output n6;
    input n30999;
    output n12138;
    input n31050;
    output n11987;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire clk_255kHz;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n2550;
    wire [31:0]n134;
    
    wire n6709, n27967, n27966, n27965, n27964, n27963, n27962, 
        n27961, n27960, n27959, n27958, n27957, n27956, n27955, 
        n27954, n27953, n27582, n27581, n27580, n27579, n27578, 
        n27577, n27576, n27575, n27574, n27573, n27572, n27571, 
        n27570, n27569, n27568, n27567, n27826, n27825, n27824, 
        n27823, n27822, n27821, n27820, n27819, n27818, n27817, 
        n27816, n27815, n27814, n27813, n27812, n27811;
    
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=508, LSE_RLINE=511 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_250 (.A(n34347), .B(clk_255kHz), .C(n6674), .Z(n32375)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_3_lut_rep_250.init = 16'h1010;
    LUT4 i24813_2_lut_rep_249_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), 
         .D(n31079), .Z(n32374)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24813_2_lut_rep_249_4_lut.init = 16'h1000;
    LUT4 i24676_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n30942), 
         .Z(n12030)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24676_2_lut_4_lut.init = 16'h1000;
    LUT4 i24759_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n31025), 
         .Z(n12031)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24759_2_lut_4_lut.init = 16'h1000;
    LUT4 i24692_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n30958), 
         .Z(n28331)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24692_2_lut_4_lut.init = 16'h1000;
    LUT4 i24674_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n30940), 
         .Z(n28339)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24674_2_lut_4_lut.init = 16'h1000;
    LUT4 i24767_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n31033), 
         .Z(n28345)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24767_2_lut_4_lut.init = 16'h1000;
    LUT4 i24775_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n31041), 
         .Z(n28337)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24775_2_lut_4_lut.init = 16'h1000;
    LUT4 i24791_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n31057), 
         .Z(n28352)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24791_2_lut_4_lut.init = 16'h1000;
    LUT4 i2_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n988), 
         .Z(n6)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_2_lut_4_lut.init = 16'h1000;
    LUT4 i24733_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n30999), 
         .Z(n12138)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24733_2_lut_4_lut.init = 16'h1000;
    LUT4 i24784_2_lut_4_lut (.A(n34347), .B(clk_255kHz), .C(n6674), .D(n31050), 
         .Z(n11987)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24784_2_lut_4_lut.init = 16'h1000;
    FD1S3IX count_2174__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2550), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i0.GSR = "ENABLED";
    FD1S3IX count_2174__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2550), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i1.GSR = "ENABLED";
    FD1S3IX count_2174__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2550), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i2.GSR = "ENABLED";
    FD1S3IX count_2174__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2550), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i3.GSR = "ENABLED";
    FD1S3IX count_2174__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2550), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i4.GSR = "ENABLED";
    FD1S3IX count_2174__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2550), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i5.GSR = "ENABLED";
    FD1S3IX count_2174__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2550), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i6.GSR = "ENABLED";
    FD1S3IX count_2174__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2550), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i7.GSR = "ENABLED";
    FD1S3IX count_2174__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2550), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i8.GSR = "ENABLED";
    FD1S3IX count_2174__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2550), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i9.GSR = "ENABLED";
    FD1S3IX count_2174__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i10.GSR = "ENABLED";
    FD1S3IX count_2174__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i11.GSR = "ENABLED";
    FD1S3IX count_2174__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i12.GSR = "ENABLED";
    FD1S3IX count_2174__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i13.GSR = "ENABLED";
    FD1S3IX count_2174__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i14.GSR = "ENABLED";
    FD1S3IX count_2174__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i15.GSR = "ENABLED";
    FD1S3IX count_2174__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i16.GSR = "ENABLED";
    FD1S3IX count_2174__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i17.GSR = "ENABLED";
    FD1S3IX count_2174__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i18.GSR = "ENABLED";
    FD1S3IX count_2174__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i19.GSR = "ENABLED";
    FD1S3IX count_2174__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i20.GSR = "ENABLED";
    FD1S3IX count_2174__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i21.GSR = "ENABLED";
    FD1S3IX count_2174__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i22.GSR = "ENABLED";
    FD1S3IX count_2174__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i23.GSR = "ENABLED";
    FD1S3IX count_2174__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i24.GSR = "ENABLED";
    FD1S3IX count_2174__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i25.GSR = "ENABLED";
    FD1S3IX count_2174__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i26.GSR = "ENABLED";
    FD1S3IX count_2174__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i27.GSR = "ENABLED";
    FD1S3IX count_2174__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i28.GSR = "ENABLED";
    FD1S3IX count_2174__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i29.GSR = "ENABLED";
    FD1S3IX count_2174__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i30.GSR = "ENABLED";
    FD1S3IX count_2174__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i31.GSR = "ENABLED";
    LUT4 i893_2_lut (.A(n6709), .B(n34347), .Z(n2550)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i893_2_lut.init = 16'heeee;
    CCU2D add_21614_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27967), 
          .S1(n6674));
    defparam add_21614_32.INIT0 = 16'h5555;
    defparam add_21614_32.INIT1 = 16'h0000;
    defparam add_21614_32.INJECT1_0 = "NO";
    defparam add_21614_32.INJECT1_1 = "NO";
    CCU2D add_21614_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27966), .COUT(n27967));
    defparam add_21614_30.INIT0 = 16'h5555;
    defparam add_21614_30.INIT1 = 16'h5555;
    defparam add_21614_30.INJECT1_0 = "NO";
    defparam add_21614_30.INJECT1_1 = "NO";
    CCU2D add_21614_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27965), .COUT(n27966));
    defparam add_21614_28.INIT0 = 16'h5555;
    defparam add_21614_28.INIT1 = 16'h5555;
    defparam add_21614_28.INJECT1_0 = "NO";
    defparam add_21614_28.INJECT1_1 = "NO";
    CCU2D add_21614_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27964), .COUT(n27965));
    defparam add_21614_26.INIT0 = 16'h5555;
    defparam add_21614_26.INIT1 = 16'h5555;
    defparam add_21614_26.INJECT1_0 = "NO";
    defparam add_21614_26.INJECT1_1 = "NO";
    CCU2D add_21614_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27963), .COUT(n27964));
    defparam add_21614_24.INIT0 = 16'h5555;
    defparam add_21614_24.INIT1 = 16'h5555;
    defparam add_21614_24.INJECT1_0 = "NO";
    defparam add_21614_24.INJECT1_1 = "NO";
    CCU2D add_21614_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27962), .COUT(n27963));
    defparam add_21614_22.INIT0 = 16'h5555;
    defparam add_21614_22.INIT1 = 16'h5555;
    defparam add_21614_22.INJECT1_0 = "NO";
    defparam add_21614_22.INJECT1_1 = "NO";
    CCU2D add_21614_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27961), .COUT(n27962));
    defparam add_21614_20.INIT0 = 16'h5555;
    defparam add_21614_20.INIT1 = 16'h5555;
    defparam add_21614_20.INJECT1_0 = "NO";
    defparam add_21614_20.INJECT1_1 = "NO";
    CCU2D add_21614_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27960), .COUT(n27961));
    defparam add_21614_18.INIT0 = 16'h5555;
    defparam add_21614_18.INIT1 = 16'h5555;
    defparam add_21614_18.INJECT1_0 = "NO";
    defparam add_21614_18.INJECT1_1 = "NO";
    CCU2D add_21614_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27959), .COUT(n27960));
    defparam add_21614_16.INIT0 = 16'h5555;
    defparam add_21614_16.INIT1 = 16'h5555;
    defparam add_21614_16.INJECT1_0 = "NO";
    defparam add_21614_16.INJECT1_1 = "NO";
    CCU2D add_21614_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27958), .COUT(n27959));
    defparam add_21614_14.INIT0 = 16'h5555;
    defparam add_21614_14.INIT1 = 16'h5555;
    defparam add_21614_14.INJECT1_0 = "NO";
    defparam add_21614_14.INJECT1_1 = "NO";
    CCU2D add_21614_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27957), .COUT(n27958));
    defparam add_21614_12.INIT0 = 16'h5555;
    defparam add_21614_12.INIT1 = 16'h5555;
    defparam add_21614_12.INJECT1_0 = "NO";
    defparam add_21614_12.INJECT1_1 = "NO";
    CCU2D add_21614_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27956), .COUT(n27957));
    defparam add_21614_10.INIT0 = 16'h5555;
    defparam add_21614_10.INIT1 = 16'h5555;
    defparam add_21614_10.INJECT1_0 = "NO";
    defparam add_21614_10.INJECT1_1 = "NO";
    CCU2D add_21614_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27955), 
          .COUT(n27956));
    defparam add_21614_8.INIT0 = 16'h5555;
    defparam add_21614_8.INIT1 = 16'h5555;
    defparam add_21614_8.INJECT1_0 = "NO";
    defparam add_21614_8.INJECT1_1 = "NO";
    CCU2D add_21614_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27954), 
          .COUT(n27955));
    defparam add_21614_6.INIT0 = 16'h5555;
    defparam add_21614_6.INIT1 = 16'h5555;
    defparam add_21614_6.INJECT1_0 = "NO";
    defparam add_21614_6.INJECT1_1 = "NO";
    CCU2D add_21614_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27953), 
          .COUT(n27954));
    defparam add_21614_4.INIT0 = 16'h5555;
    defparam add_21614_4.INIT1 = 16'h5aaa;
    defparam add_21614_4.INJECT1_0 = "NO";
    defparam add_21614_4.INJECT1_1 = "NO";
    CCU2D add_21614_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27953));
    defparam add_21614_2.INIT0 = 16'h7000;
    defparam add_21614_2.INIT1 = 16'h5aaa;
    defparam add_21614_2.INJECT1_0 = "NO";
    defparam add_21614_2.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27582), .S0(n6709));
    defparam sub_1709_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1709_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1709_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1709_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27581), .COUT(n27582));
    defparam sub_1709_add_2_32.INIT0 = 16'h5555;
    defparam sub_1709_add_2_32.INIT1 = 16'h5555;
    defparam sub_1709_add_2_32.INJECT1_0 = "NO";
    defparam sub_1709_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27580), .COUT(n27581));
    defparam sub_1709_add_2_30.INIT0 = 16'h5555;
    defparam sub_1709_add_2_30.INIT1 = 16'h5555;
    defparam sub_1709_add_2_30.INJECT1_0 = "NO";
    defparam sub_1709_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27579), .COUT(n27580));
    defparam sub_1709_add_2_28.INIT0 = 16'h5555;
    defparam sub_1709_add_2_28.INIT1 = 16'h5555;
    defparam sub_1709_add_2_28.INJECT1_0 = "NO";
    defparam sub_1709_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27578), .COUT(n27579));
    defparam sub_1709_add_2_26.INIT0 = 16'h5555;
    defparam sub_1709_add_2_26.INIT1 = 16'h5555;
    defparam sub_1709_add_2_26.INJECT1_0 = "NO";
    defparam sub_1709_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27577), .COUT(n27578));
    defparam sub_1709_add_2_24.INIT0 = 16'h5555;
    defparam sub_1709_add_2_24.INIT1 = 16'h5555;
    defparam sub_1709_add_2_24.INJECT1_0 = "NO";
    defparam sub_1709_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27576), .COUT(n27577));
    defparam sub_1709_add_2_22.INIT0 = 16'h5555;
    defparam sub_1709_add_2_22.INIT1 = 16'h5555;
    defparam sub_1709_add_2_22.INJECT1_0 = "NO";
    defparam sub_1709_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27575), .COUT(n27576));
    defparam sub_1709_add_2_20.INIT0 = 16'h5555;
    defparam sub_1709_add_2_20.INIT1 = 16'h5555;
    defparam sub_1709_add_2_20.INJECT1_0 = "NO";
    defparam sub_1709_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27574), .COUT(n27575));
    defparam sub_1709_add_2_18.INIT0 = 16'h5555;
    defparam sub_1709_add_2_18.INIT1 = 16'h5555;
    defparam sub_1709_add_2_18.INJECT1_0 = "NO";
    defparam sub_1709_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27573), .COUT(n27574));
    defparam sub_1709_add_2_16.INIT0 = 16'h5555;
    defparam sub_1709_add_2_16.INIT1 = 16'h5555;
    defparam sub_1709_add_2_16.INJECT1_0 = "NO";
    defparam sub_1709_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27572), .COUT(n27573));
    defparam sub_1709_add_2_14.INIT0 = 16'h5555;
    defparam sub_1709_add_2_14.INIT1 = 16'h5555;
    defparam sub_1709_add_2_14.INJECT1_0 = "NO";
    defparam sub_1709_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27571), .COUT(n27572));
    defparam sub_1709_add_2_12.INIT0 = 16'h5555;
    defparam sub_1709_add_2_12.INIT1 = 16'h5555;
    defparam sub_1709_add_2_12.INJECT1_0 = "NO";
    defparam sub_1709_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27570), .COUT(n27571));
    defparam sub_1709_add_2_10.INIT0 = 16'h5555;
    defparam sub_1709_add_2_10.INIT1 = 16'h5555;
    defparam sub_1709_add_2_10.INJECT1_0 = "NO";
    defparam sub_1709_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27569), .COUT(n27570));
    defparam sub_1709_add_2_8.INIT0 = 16'h5555;
    defparam sub_1709_add_2_8.INIT1 = 16'h5555;
    defparam sub_1709_add_2_8.INJECT1_0 = "NO";
    defparam sub_1709_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27568), .COUT(n27569));
    defparam sub_1709_add_2_6.INIT0 = 16'h5555;
    defparam sub_1709_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_1709_add_2_6.INJECT1_0 = "NO";
    defparam sub_1709_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27567), .COUT(n27568));
    defparam sub_1709_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1709_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_1709_add_2_4.INJECT1_0 = "NO";
    defparam sub_1709_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27567));
    defparam sub_1709_add_2_2.INIT0 = 16'h0000;
    defparam sub_1709_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1709_add_2_2.INJECT1_0 = "NO";
    defparam sub_1709_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27826), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_33.INIT1 = 16'h0000;
    defparam count_2174_add_4_33.INJECT1_0 = "NO";
    defparam count_2174_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27825), .COUT(n27826), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_31.INJECT1_0 = "NO";
    defparam count_2174_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27824), .COUT(n27825), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_29.INJECT1_0 = "NO";
    defparam count_2174_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27823), .COUT(n27824), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_27.INJECT1_0 = "NO";
    defparam count_2174_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27822), .COUT(n27823), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_25.INJECT1_0 = "NO";
    defparam count_2174_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27821), .COUT(n27822), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_23.INJECT1_0 = "NO";
    defparam count_2174_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27820), .COUT(n27821), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_21.INJECT1_0 = "NO";
    defparam count_2174_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27819), .COUT(n27820), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_19.INJECT1_0 = "NO";
    defparam count_2174_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27818), .COUT(n27819), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_17.INJECT1_0 = "NO";
    defparam count_2174_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27817), .COUT(n27818), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_15.INJECT1_0 = "NO";
    defparam count_2174_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27816), .COUT(n27817), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_13.INJECT1_0 = "NO";
    defparam count_2174_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27815), .COUT(n27816), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_11.INJECT1_0 = "NO";
    defparam count_2174_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27814), .COUT(n27815), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_9.INJECT1_0 = "NO";
    defparam count_2174_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27813), .COUT(n27814), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_7.INJECT1_0 = "NO";
    defparam count_2174_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27812), .COUT(n27813), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_5.INJECT1_0 = "NO";
    defparam count_2174_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27811), .COUT(n27812), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_3.INJECT1_0 = "NO";
    defparam count_2174_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27811), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_1.INIT0 = 16'hF000;
    defparam count_2174_add_4_1.INIT1 = 16'h0555;
    defparam count_2174_add_4_1.INJECT1_0 = "NO";
    defparam count_2174_add_4_1.INJECT1_1 = "NO";
    
endmodule
