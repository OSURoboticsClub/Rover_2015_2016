// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Mon Apr 25 18:00:08 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(362[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    inout expansion4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[13:23])
    input expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire n33383 /* synthesis nomerge= */ ;
    
    wire GND_net, VCC_net, uart_rx_c, n11072, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, expansion1_c_9, expansion2_c_10, expansion3_c_11, 
        expansion5_c, signal_light_c, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
        encoder_la_c, encoder_lb_c, encoder_li_c, rc_ch1_c, rc_ch2_c, 
        rc_ch3_c, rc_ch4_c, rc_ch7_c, rc_ch8_c, motor_pwm_l_c, xbee_pause_c, 
        debug_c_7, debug_c_5, debug_c_4, debug_c_3, debug_c_2, debug_c_0;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(451[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(452[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    
    wire rw, n14453, n14546;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    
    wire timeout_pause;
    wire [31:0]timeout_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[13:26])
    
    wire prev_uart_rx, clk_255kHz, n27751, n27549, n14650, n1155, 
        n8, n9, n2;
    wire [31:0]n99_adj_1336;
    wire [7:0]n8634;
    
    wire n2_adj_605;
    wire [31:0]n100_adj_1355;
    wire [31:0]n657;
    
    wire n35;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n21208, n13, n21211, n14, n21213, n6, n15086, n2966, 
        n21219, n21221;
    wire [31:0]n1473;
    
    wire n12, n29901, n29256, n14522, n31445, n29826, n5833, n8506, 
        n9368, n2875, n2869, n14513, n14512, n3, n2_adj_606, n27444;
    wire [31:0]n5973;
    
    wire n29943, n2860, n2857, n10, n32, n13315, n3_adj_607, n8_adj_608, 
        n24, n2_adj_609, n9537, n4006, force_pause;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    
    wire clk_1Hz, prev_clk_1Hz;
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(32[12:21])
    
    wire n46, n22395, n22389, n14145, n31409;
    wire [7:0]\register[0]_adj_975 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]read_value_adj_976;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(92[12:22])
    
    wire n22;
    wire [2:0]read_size_adj_977;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(93[12:21])
    
    wire n64, n32_adj_619, n16842, n16841, n34, n27535, n29236, 
        n3_adj_620, n27441, n2846, n14499, n16840, n241, n27427, 
        n9330;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched, prev_limit_latched, step_clk, prev_step_clk;
    wire [31:0]read_value_adj_983;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_984;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select, n52, n17, n16, n15, n303, n31444, n31443, 
        n73, n18, n16012, n4180;
    wire [7:0]control_reg_adj_992;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_993;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_994;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched_adj_656, prev_limit_latched_adj_657, int_step, 
        step_clk_adj_658, prev_step_clk_adj_659;
    wire [31:0]read_value_adj_995;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_996;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_694, n4, n52_adj_695;
    wire [31:0]n224_adj_999;
    
    wire n27168, n27167, n27166, n27165, n8401, n31442, n27164;
    wire [31:0]n4094;
    
    wire n27163, n27162, n8_adj_697, n8367, n14_adj_698, n13_adj_699, 
        n27161, n27160, n2_adj_700, n33387, n27159, n27158, n3_adj_701;
    wire [31:0]steps_reg_adj_1033;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched_adj_702, prev_limit_latched_adj_703;
    wire [31:0]read_value_adj_1034;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_1035;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_738, n8_adj_739, n11, n8_adj_740, n2_adj_741, 
        n13956, n9304, n13947, n2_adj_742, n8055, n13940, n33386;
    wire [31:0]n580_adj_1053;
    
    wire n13938, n9300, n5;
    wire [7:0]control_reg_adj_1070;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched_adj_744, prev_limit_latched_adj_745;
    wire [31:0]read_value_adj_1073;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_1074;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_780, n29837;
    wire [31:0]n224_adj_1077;
    
    wire n8297, n8_adj_813, n31410, n8_adj_814, n8_adj_815;
    wire [31:0]n3921;
    
    wire n27542, n13916, n2_adj_816, n9483, n29783, n9296, n29491, 
        n13907, n2_adj_817, n8263, n8_adj_818, n31408, n2823;
    wire [31:0]\register[1]_adj_1109 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    wire qreset;
    wire [31:0]read_value_adj_1111;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(65[13:23])
    wire [2:0]read_size_adj_1112;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[12:21])
    
    wire prev_select_adj_853;
    wire [31:0]read_value_adj_1119;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(65[13:23])
    wire [2:0]read_size_adj_1120;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[12:21])
    
    wire prev_select_adj_888;
    wire [7:0]\register[1]_adj_1133 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]\register[0]_adj_1134 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]read_value_adj_1135;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(26[12:22])
    wire [2:0]read_size_adj_1136;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(27[12:21])
    
    wire prev_select_adj_898, n176, n31412, n13833, n29234, n29293, 
        n29300, n9_adj_899, n29292, n2_adj_900, n3_adj_901, n2_adj_902, 
        n2_adj_903, n8_adj_904;
    wire [14:0]n33690;
    
    wire n8_adj_906, n12210, n31411, n31435, n31434, n31431, n31427, 
        n31426, n31425, n31424, n6_adj_907, n33384, n27679, n29817, 
        n1, n2_adj_908, n8_adj_909, n14_adj_910, n2_adj_911, n2_adj_912, 
        n8_adj_913, n24145, n29791, n2_adj_914, n29846, n2_adj_915, 
        n8_adj_916, n2_adj_917, n2_adj_918, n8_adj_919, n8_adj_920, 
        n29810, n2_adj_921, n8_adj_922, n2_adj_923, n8_adj_924, n29788, 
        n2_adj_925, n2_adj_926, n12148, n8_adj_927, n8_adj_928, n2_adj_929, 
        n2_adj_930, n8_adj_931, n3_adj_932, n2_adj_933, n2_adj_934, 
        n8_adj_935, n29169, n2_adj_936, n29529, n26434, n29839;
    wire [7:0]n8652;
    
    wire n56, n26433, n66, n2_adj_937, n22483, n9_adj_938, n8193, 
        n26432, n14782, n31600, n27540, n11235;
    wire [31:0]n6778;
    
    wire n30, n26431, n26430, n31595, n17034, select_clk, n9378, 
        n26429, n31590, n31589, n26428, n26427, n26426, n31587, 
        n31421, n26425;
    wire [1:0]n33623;
    
    wire n31581, n42, n40, n38, n36, n34_adj_940, expansion4_out, 
        n31575, n30_adj_941, n29, n30305, n26, n29270, n31570, 
        n26424, n29136, n31555, n11007, n33385, n11208, n2_adj_942, 
        n2_adj_943, n29263, n6_adj_944, n12368, n31540, n31539, 
        n29333, n31536, n7916, n21502, n31532, n27563;
    wire [2:0]quadA_delayed_adj_1223;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [2:0]quadB_delayed_adj_1224;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n31529, n8159, n33389, n27752, n8_adj_945, n8_adj_946, 
        n29113, n11006, n31525, n12158, n9580, n9547, n9541, n3_adj_947, 
        n30303, n31511, n7881, n29199, n29066, n28826, n29056, 
        n29053, n29065, n29063, n29050, n29052, n29054, n31503, 
        n29067, n29057, n31501, n27546, n29068, n29071, n31500, 
        n29070, n27464, n31496, n29058, n29059, n29064, n29060, 
        n29062, n31406, n29055, n29051, n31407, n29049, n29061, 
        n29048, n29069, n29294, n29220, n3_adj_948, n31420, n29831, 
        n7846, n27483, n8089, n29257, n31482, n29112, n27249, 
        n31477, n31476, n31473, n31472, n31419, n31470, n31469, 
        n31465, n16764, n31464, n29331, n31463, n31418, n31462, 
        n26423, n26422, n26421, n26420, n31456, n26419, n107;
    wire [3:0]state_adj_1312;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n29047, n26889, n26888, n13155, n27784, n31449, n26887, 
        n26886, n29829, n26885, n26884, n31448, n26883, n16763, 
        n31446, n29785;
    
    VHI i2 (.Z(VCC_net));
    ExpansionGPIO gpio (.read_value({read_value_adj_1135}), .debug_c_c(debug_c_c), 
            .n2869(n2869), .n29220(n29220), .n13947(n13947), .n31511(n31511), 
            .\databus[0] (databus[0]), .\read_size[0] (read_size_adj_1136[0]), 
            .n27679(n27679), .prev_select(prev_select_adj_898), .\select[5] (select[5]), 
            .expansion1_c_9(expansion1_c_9), .n31435(n31435), .n56(n56), 
            .expansion2_c_10(expansion2_c_10), .expansion3_c_11(expansion3_c_11), 
            .\databus[1] (databus[1]), .\databus[2] (databus[2]), .\databus[3] (databus[3]), 
            .\register[0][4] (\register[0]_adj_1134 [4]), .\databus[4] (databus[4]), 
            .\register[0][5] (\register[0]_adj_1134 [5]), .\databus[5] (databus[5]), 
            .\databus[6] (databus[6]), .\databus[7] (databus[7]), .n16012(n16012), 
            .\register[1][4] (\register[1]_adj_1133 [4]), .\register[1][5] (\register[1]_adj_1133 [5]), 
            .n12368(n12368), .n31406(n31406), .\register_addr[0] (register_addr[0]), 
            .n24145(n24145), .n11007(n11007), .n11006(n11006)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(692[18] 703[38])
    IFS1P3DX prev_uart_rx_57 (.D(uart_rx_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(prev_uart_rx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam prev_uart_rx_57.GSR = "ENABLED";
    FD1S3AX timeout_pause_59 (.D(n27784), .CK(debug_c_c), .Q(timeout_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_pause_59.GSR = "ENABLED";
    LUT4 i1043_2_lut_rep_266_3_lut (.A(n22483), .B(reset_count[14]), .C(n8367), 
         .Z(n31409)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1043_2_lut_rep_266_3_lut.init = 16'hf7f7;
    LUT4 i15031_2_lut_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(databus[4]), 
         .Z(n580_adj_1053[4])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15031_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_rep_269_4_lut (.A(n22483), .B(reset_count[14]), .C(n8506), 
         .D(select_clk), .Z(n31412)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_269_4_lut.init = 16'h0080;
    CCU2D add_30_9 (.A0(timeout_count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26422), .COUT(n26423), .S0(n657[7]), .S1(n657[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_9.INIT0 = 16'h5aaa;
    defparam add_30_9.INIT1 = 16'h5aaa;
    defparam add_30_9.INJECT1_0 = "NO";
    defparam add_30_9.INJECT1_1 = "NO";
    CCU2D add_30_7 (.A0(timeout_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26421), .COUT(n26422), .S0(n657[5]), .S1(n657[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_7.INIT0 = 16'h5aaa;
    defparam add_30_7.INIT1 = 16'h5aaa;
    defparam add_30_7.INJECT1_0 = "NO";
    defparam add_30_7.INJECT1_1 = "NO";
    LUT4 i10291_2_lut_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(n8089), 
         .D(n8055), .Z(n17034)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10291_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i14814_2_lut_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(n7881), 
         .Z(n241)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i14814_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i5444_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(limit_latched_adj_744), 
         .D(prev_limit_latched_adj_745), .Z(n12210)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i5444_3_lut_4_lut.init = 16'h77f7;
    LUT4 i22481_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(n73), 
         .D(state_adj_1312[2]), .Z(n14782)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i22481_3_lut_4_lut.init = 16'hff7f;
    LUT4 i22344_4_lut (.A(n29333), .B(reset_count[14]), .C(n13315), .D(n21502), 
         .Z(n30)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i22344_4_lut.init = 16'h373f;
    LUT4 i1_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(n9304), .Z(n14546)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut (.A(n22395), .B(n29331), .C(reset_count[6]), .D(reset_count[5]), 
         .Z(n29333)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(461[7:30])
    defparam i1_4_lut.init = 16'hfcec;
    LUT4 i1_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(prev_limit_latched_adj_703), 
         .D(limit_latched_adj_702), .Z(n11208)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h7f77;
    LUT4 i15652_4_lut (.A(reset_count[0]), .B(reset_count[4]), .C(n6_adj_907), 
         .D(reset_count[3]), .Z(n22395)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i15652_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(reset_count[1]), .B(reset_count[2]), .Z(n6_adj_907)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(reset_count[11]), .B(reset_count[12]), .C(reset_count[13]), 
         .Z(n13315)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(461[7:30])
    defparam i2_3_lut.init = 16'hfefe;
    VLO i1 (.Z(GND_net));
    LUT4 i4_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(debug_c_0), 
         .Z(qreset)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i4_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_3_lut_4_lut_adj_509 (.A(n22483), .B(reset_count[14]), .C(prev_limit_latched), 
         .D(limit_latched), .Z(n12158)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_509.init = 16'h7f77;
    LUT4 i5383_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(limit_latched_adj_656), 
         .D(prev_limit_latched_adj_657), .Z(n12148)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i5383_3_lut_4_lut.init = 16'h77f7;
    LUT4 i22327_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(n29785), 
         .Z(n2966)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i22327_2_lut_3_lut.init = 16'hf7f7;
    FD1P3IX timeout_count__i0 (.D(n100_adj_1355[0]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i0.GSR = "ENABLED";
    LUT4 i22330_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(n29788), 
         .Z(n2875)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i22330_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i22333_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(n29791), 
         .Z(n2860)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i22333_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i973_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(n7916), 
         .Z(n2823)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i973_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1031_2_lut_rep_265_3_lut (.A(n22483), .B(reset_count[14]), .C(n8055), 
         .Z(n31408)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1031_2_lut_rep_265_3_lut.init = 16'hf7f7;
    LUT4 i10068_2_lut_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(n8193), 
         .D(n8159), .Z(n16840)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10068_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1035_2_lut_rep_264_3_lut (.A(n22483), .B(reset_count[14]), .C(n8159), 
         .Z(n31407)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1035_2_lut_rep_264_3_lut.init = 16'hf7f7;
    CCU2D add_30_5 (.A0(timeout_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26420), .COUT(n26421), .S0(n100_adj_1355[3]), 
          .S1(n657[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_5.INIT0 = 16'h5aaa;
    defparam add_30_5.INIT1 = 16'h5aaa;
    defparam add_30_5.INJECT1_0 = "NO";
    defparam add_30_5.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_268_4_lut (.A(n22483), .B(reset_count[14]), .C(n7881), 
         .D(clk_255kHz), .Z(n31411)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_268_4_lut.init = 16'h0080;
    LUT4 i1_3_lut_rep_319_4_lut (.A(n22483), .B(reset_count[14]), .C(state_adj_1312[3]), 
         .D(state_adj_1312[2]), .Z(n31462)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_319_4_lut.init = 16'h0888;
    LUT4 i2758_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(prev_clk_1Hz), 
         .D(clk_1Hz), .Z(n9483)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i2758_3_lut_4_lut.init = 16'h7f77;
    LUT4 i10069_2_lut_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(n8297), 
         .D(n8263), .Z(n16841)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10069_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1039_2_lut_rep_267_3_lut (.A(n22483), .B(reset_count[14]), .C(n8263), 
         .Z(n31410)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1039_2_lut_rep_267_3_lut.init = 16'hf7f7;
    LUT4 i15229_2_lut_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(n8506), 
         .Z(n107)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15229_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i10070_2_lut_3_lut_4_lut (.A(n22483), .B(reset_count[14]), .C(n8401), 
         .D(n8367), .Z(n16842)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10070_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i14850_2_lut_2_lut_3_lut (.A(n22483), .B(reset_count[14]), .C(databus[2]), 
         .Z(n580_adj_1053[2])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i14850_2_lut_2_lut_3_lut.init = 16'h8080;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i2_3_lut_rep_288_4_lut (.A(select[3]), .B(n31501), .C(n31525), 
         .D(prev_select_adj_888), .Z(n31431)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam i2_3_lut_rep_288_4_lut.init = 16'h0080;
    LUT4 Select_4295_i10_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1119[1]), 
         .D(n33384), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4295_i10_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_3_lut (.A(n31500), .B(n1473[17]), .C(n1473[20]), .Z(n27464)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i2_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i22362_4_lut_4_lut (.A(n31500), .B(n4), .C(n5833), .D(n1473[14]), 
         .Z(n13833)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i22362_4_lut_4_lut.init = 16'h2a00;
    LUT4 i2_3_lut_rep_469 (.A(n22483), .B(reset_count[14]), .C(n7881), 
         .D(clk_255kHz), .Z(n33387)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_469.init = 16'h0080;
    CCU2D add_19622_24 (.A0(timeout_count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27168), .S1(n7846));
    defparam add_19622_24.INIT0 = 16'h5555;
    defparam add_19622_24.INIT1 = 16'h0000;
    defparam add_19622_24.INJECT1_0 = "NO";
    defparam add_19622_24.INJECT1_1 = "NO";
    CCU2D add_19622_22 (.A0(timeout_count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27167), .COUT(n27168));
    defparam add_19622_22.INIT0 = 16'h5555;
    defparam add_19622_22.INIT1 = 16'h5555;
    defparam add_19622_22.INJECT1_0 = "NO";
    defparam add_19622_22.INJECT1_1 = "NO";
    CCU2D add_19622_20 (.A0(timeout_count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27166), .COUT(n27167));
    defparam add_19622_20.INIT0 = 16'h5555;
    defparam add_19622_20.INIT1 = 16'h5555;
    defparam add_19622_20.INJECT1_0 = "NO";
    defparam add_19622_20.INJECT1_1 = "NO";
    CCU2D add_19622_18 (.A0(timeout_count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27165), .COUT(n27166));
    defparam add_19622_18.INIT0 = 16'h5aaa;
    defparam add_19622_18.INIT1 = 16'h5555;
    defparam add_19622_18.INJECT1_0 = "NO";
    defparam add_19622_18.INJECT1_1 = "NO";
    CCU2D add_19622_16 (.A0(timeout_count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27164), .COUT(n27165));
    defparam add_19622_16.INIT0 = 16'h5aaa;
    defparam add_19622_16.INIT1 = 16'h5aaa;
    defparam add_19622_16.INJECT1_0 = "NO";
    defparam add_19622_16.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n31511), .B(prev_select_adj_780), 
         .C(n31465), .D(register_addr[5]), .Z(n2857)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    CCU2D add_19622_14 (.A0(timeout_count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27163), .COUT(n27164));
    defparam add_19622_14.INIT0 = 16'h5555;
    defparam add_19622_14.INIT1 = 16'h5555;
    defparam add_19622_14.INJECT1_0 = "NO";
    defparam add_19622_14.INJECT1_1 = "NO";
    CCU2D add_19622_12 (.A0(timeout_count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27162), .COUT(n27163));
    defparam add_19622_12.INIT0 = 16'h5555;
    defparam add_19622_12.INIT1 = 16'h5aaa;
    defparam add_19622_12.INJECT1_0 = "NO";
    defparam add_19622_12.INJECT1_1 = "NO";
    CCU2D add_19622_10 (.A0(timeout_count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27161), .COUT(n27162));
    defparam add_19622_10.INIT0 = 16'h5aaa;
    defparam add_19622_10.INIT1 = 16'h5555;
    defparam add_19622_10.INJECT1_0 = "NO";
    defparam add_19622_10.INJECT1_1 = "NO";
    CCU2D add_19622_8 (.A0(timeout_count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27160), .COUT(n27161));
    defparam add_19622_8.INIT0 = 16'h5aaa;
    defparam add_19622_8.INIT1 = 16'h5aaa;
    defparam add_19622_8.INJECT1_0 = "NO";
    defparam add_19622_8.INJECT1_1 = "NO";
    CCU2D add_19622_6 (.A0(timeout_count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27159), .COUT(n27160));
    defparam add_19622_6.INIT0 = 16'h5555;
    defparam add_19622_6.INIT1 = 16'h5555;
    defparam add_19622_6.INJECT1_0 = "NO";
    defparam add_19622_6.INJECT1_1 = "NO";
    CCU2D add_19622_4 (.A0(timeout_count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27158), .COUT(n27159));
    defparam add_19622_4.INIT0 = 16'h5555;
    defparam add_19622_4.INIT1 = 16'h5555;
    defparam add_19622_4.INJECT1_0 = "NO";
    defparam add_19622_4.INJECT1_1 = "NO";
    LUT4 i22442_4_lut (.A(n29901), .B(n17), .C(n15), .D(n16), .Z(n27784)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i22442_4_lut.init = 16'h8000;
    CCU2D add_19622_2 (.A0(timeout_count[9]), .B0(timeout_count[8]), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27158));
    defparam add_19622_2.INIT0 = 16'h7000;
    defparam add_19622_2.INIT1 = 16'h5aaa;
    defparam add_19622_2.INJECT1_0 = "NO";
    defparam add_19622_2.INJECT1_1 = "NO";
    LUT4 i22441_4_lut (.A(n29), .B(n42), .C(n38), .D(n30_adj_941), .Z(n29901)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i22441_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(timeout_count[16]), .B(timeout_count[25]), .C(timeout_count[15]), 
         .D(timeout_count[24]), .Z(n17)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(timeout_count[8]), .B(timeout_count[20]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i6_4_lut (.A(timeout_count[17]), .B(timeout_count[9]), .C(timeout_count[23]), 
         .D(timeout_count[10]), .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i7_2_lut (.A(timeout_count[5]), .B(timeout_count[18]), .Z(n29)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(timeout_count[12]), .B(n40), .C(n34_adj_940), .D(timeout_count[19]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(timeout_count[31]), .B(timeout_count[22]), .C(timeout_count[21]), 
         .D(timeout_count[28]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i16_4_lut.init = 16'hfffe;
    FD1P3AX reset_count_2668_2669__i1 (.D(n33690[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i1.GSR = "ENABLED";
    LUT4 i8_2_lut (.A(timeout_count[1]), .B(timeout_count[4]), .Z(n30_adj_941)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(timeout_count[6]), .B(n36), .C(n26), .D(timeout_count[2]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i12_4_lut (.A(timeout_count[14]), .B(timeout_count[11]), .C(timeout_count[30]), 
         .D(timeout_count[13]), .Z(n34_adj_940)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(timeout_count[29]), .B(timeout_count[26]), .C(timeout_count[7]), 
         .D(timeout_count[3]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(timeout_count[0]), .B(timeout_count[27]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_rep_357 (.A(reset_count[14]), .B(reset_count[12]), .C(reset_count[13]), 
         .D(n29263), .Z(n31500)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam i1_4_lut_rep_357.init = 16'hfaea;
    LUT4 i15745_1_lut_rep_329_4_lut (.A(reset_count[14]), .B(reset_count[12]), 
         .C(reset_count[13]), .D(n29263), .Z(n31472)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam i15745_1_lut_rep_329_4_lut.init = 16'h0515;
    LUT4 i15_2_lut_rep_300_3_lut_4_lut (.A(register_addr[4]), .B(n31532), 
         .C(rw), .D(select[3]), .Z(n31443)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam i15_2_lut_rep_300_3_lut_4_lut.init = 16'hd000;
    LUT4 i114_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n31532), .C(prev_select_adj_853), 
         .D(select[3]), .Z(n14145)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam i114_2_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 Select_4300_i6_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n31532), 
         .C(read_size_adj_1112[2]), .D(select[3]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4300_i6_2_lut_3_lut_4_lut.init = 16'hd000;
    LUT4 i15_2_lut_rep_303_3_lut_4_lut (.A(register_addr[4]), .B(n31532), 
         .C(rw), .D(select[3]), .Z(n31446)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam i15_2_lut_rep_303_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4307_i9_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n31532), 
         .C(read_size_adj_1120[0]), .D(select[3]), .Z(n9)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4307_i9_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i114_2_lut_3_lut_4_lut_adj_510 (.A(register_addr[4]), .B(n31532), 
         .C(prev_select_adj_888), .D(select[3]), .Z(n15086)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam i114_2_lut_3_lut_4_lut_adj_510.init = 16'h0200;
    LUT4 i2_3_lut_rep_467 (.A(n22483), .B(reset_count[14]), .C(n7881), 
         .D(clk_255kHz), .Z(n33385)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_467.init = 16'h0080;
    LUT4 i2_3_lut_rep_468 (.A(n22483), .B(reset_count[14]), .C(n7881), 
         .D(clk_255kHz), .Z(n33386)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_468.init = 16'h0080;
    LUT4 i22420_2_lut_rep_368 (.A(n22483), .B(reset_count[14]), .Z(n31511)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22420_2_lut_rep_368.init = 16'h7777;
    CCU2D add_30_3 (.A0(timeout_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26419), .COUT(n26420), .S0(n100_adj_1355[1]), 
          .S1(n100_adj_1355[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_3.INIT0 = 16'h5aaa;
    defparam add_30_3.INIT1 = 16'h5aaa;
    defparam add_30_3.INJECT1_0 = "NO";
    defparam add_30_3.INJECT1_1 = "NO";
    LUT4 Select_4231_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[27]), 
         .D(n33384), .Z(n8_adj_814)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4231_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    CCU2D add_30_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(timeout_count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26419), .S1(n100_adj_1355[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_1.INIT0 = 16'hF000;
    defparam add_30_1.INIT1 = 16'h5555;
    defparam add_30_1.INJECT1_0 = "NO";
    defparam add_30_1.INJECT1_1 = "NO";
    LUT4 i14773_2_lut (.A(reset_count[9]), .B(reset_count[10]), .Z(n21502)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14773_2_lut.init = 16'h8888;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    IB encoder_li_pad (.I(encoder_li), .O(encoder_li_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    IB encoder_lb_pad (.I(encoder_lb), .O(encoder_lb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    IB encoder_la_pad (.I(encoder_la), .O(encoder_la_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    IB encoder_ri_pad (.I(encoder_ri), .O(encoder_ri_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    IB encoder_rb_pad (.I(encoder_rb), .O(encoder_rb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    IB encoder_ra_pad (.I(encoder_ra), .O(encoder_ra_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    IB expansion5_pad (.I(expansion5), .O(expansion5_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    IB uart_rx_pad (.I(uart_rx), .O(uart_rx_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    OB debug_pad_0 (.I(debug_c_0), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_1 (.I(n11072), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_6 (.I(n31511), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB motor_pwm_r_pad (.I(GND_net), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    OB expansion3_pad (.I(expansion3_c_11), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion2_pad (.I(expansion2_c_10), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB expansion1_pad (.I(expansion1_c_9), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    CCU2D add_30_33 (.A0(timeout_count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26434), .S0(n657[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_33.INIT0 = 16'h5aaa;
    defparam add_30_33.INIT1 = 16'h0000;
    defparam add_30_33.INJECT1_0 = "NO";
    defparam add_30_33.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_4_lut (.A(n31511), .B(n31581), .C(n31476), .D(register_addr[1]), 
         .Z(n9541)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 Select_4234_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[26]), 
         .D(n33384), .Z(n8_adj_913)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4234_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    CCU2D add_30_31 (.A0(timeout_count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26433), .COUT(n26434), .S0(n657[29]), 
          .S1(n657[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_31.INIT0 = 16'h5aaa;
    defparam add_30_31.INIT1 = 16'h5aaa;
    defparam add_30_31.INJECT1_0 = "NO";
    defparam add_30_31.INJECT1_1 = "NO";
    CCU2D add_30_17 (.A0(timeout_count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26426), .COUT(n26427), .S0(n657[15]), 
          .S1(n657[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_17.INIT0 = 16'h5aaa;
    defparam add_30_17.INIT1 = 16'h5aaa;
    defparam add_30_17.INJECT1_0 = "NO";
    defparam add_30_17.INJECT1_1 = "NO";
    CCU2D add_30_29 (.A0(timeout_count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26432), .COUT(n26433), .S0(n657[27]), 
          .S1(n657[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_29.INIT0 = 16'h5aaa;
    defparam add_30_29.INIT1 = 16'h5aaa;
    defparam add_30_29.INJECT1_0 = "NO";
    defparam add_30_29.INJECT1_1 = "NO";
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    CCU2D add_30_15 (.A0(timeout_count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26425), .COUT(n26426), .S0(n657[13]), 
          .S1(n657[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_15.INIT0 = 16'h5aaa;
    defparam add_30_15.INIT1 = 16'h5aaa;
    defparam add_30_15.INJECT1_0 = "NO";
    defparam add_30_15.INJECT1_1 = "NO";
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB uart_tx_pad (.I(n11072), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    BB expansion4_pad (.I(n11007), .T(n11006), .B(expansion4), .O(expansion4_out));
    CCU2D add_30_13 (.A0(timeout_count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26424), .COUT(n26425), .S0(n657[11]), 
          .S1(n657[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_13.INIT0 = 16'h5aaa;
    defparam add_30_13.INIT1 = 16'h5aaa;
    defparam add_30_13.INJECT1_0 = "NO";
    defparam add_30_13.INJECT1_1 = "NO";
    FD1P3IX timeout_count__i1 (.D(n100_adj_1355[1]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i1.GSR = "ENABLED";
    FD1P3IX timeout_count__i2 (.D(n100_adj_1355[2]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i2.GSR = "ENABLED";
    FD1P3IX timeout_count__i3 (.D(n100_adj_1355[3]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i3.GSR = "ENABLED";
    FD1P3IX timeout_count__i4 (.D(n657[4]), .SP(n9368), .CD(n9580), .CK(debug_c_c), 
            .Q(timeout_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i4.GSR = "ENABLED";
    FD1P3IX timeout_count__i5 (.D(n657[5]), .SP(n9368), .CD(n9580), .CK(debug_c_c), 
            .Q(timeout_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i5.GSR = "ENABLED";
    FD1P3IX timeout_count__i6 (.D(n657[6]), .SP(n9368), .CD(n9580), .CK(debug_c_c), 
            .Q(timeout_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i6.GSR = "ENABLED";
    FD1P3IX timeout_count__i7 (.D(n657[7]), .SP(n9368), .CD(n9580), .CK(debug_c_c), 
            .Q(timeout_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i7.GSR = "ENABLED";
    FD1P3IX timeout_count__i8 (.D(n657[8]), .SP(n9368), .CD(n9580), .CK(debug_c_c), 
            .Q(timeout_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i8.GSR = "ENABLED";
    FD1P3IX timeout_count__i9 (.D(n657[9]), .SP(n9368), .CD(n9580), .CK(debug_c_c), 
            .Q(timeout_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i9.GSR = "ENABLED";
    FD1P3IX timeout_count__i10 (.D(n657[10]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i10.GSR = "ENABLED";
    FD1P3IX timeout_count__i11 (.D(n657[11]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i11.GSR = "ENABLED";
    FD1P3IX timeout_count__i12 (.D(n657[12]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i12.GSR = "ENABLED";
    FD1P3IX timeout_count__i13 (.D(n657[13]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i13.GSR = "ENABLED";
    FD1P3IX timeout_count__i14 (.D(n657[14]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i14.GSR = "ENABLED";
    FD1P3IX timeout_count__i15 (.D(n657[15]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i15.GSR = "ENABLED";
    FD1P3IX timeout_count__i16 (.D(n657[16]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i16.GSR = "ENABLED";
    FD1P3IX timeout_count__i17 (.D(n657[17]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i17.GSR = "ENABLED";
    FD1P3IX timeout_count__i18 (.D(n657[18]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i18.GSR = "ENABLED";
    FD1P3IX timeout_count__i19 (.D(n657[19]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i19.GSR = "ENABLED";
    FD1P3IX timeout_count__i20 (.D(n657[20]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i20.GSR = "ENABLED";
    FD1P3IX timeout_count__i21 (.D(n657[21]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i21.GSR = "ENABLED";
    FD1P3IX timeout_count__i22 (.D(n657[22]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i22.GSR = "ENABLED";
    FD1P3IX timeout_count__i23 (.D(n657[23]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i23.GSR = "ENABLED";
    FD1P3IX timeout_count__i24 (.D(n657[24]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i24.GSR = "ENABLED";
    FD1P3IX timeout_count__i25 (.D(n657[25]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i25.GSR = "ENABLED";
    FD1P3IX timeout_count__i26 (.D(n657[26]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i26.GSR = "ENABLED";
    FD1P3IX timeout_count__i27 (.D(n657[27]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i27.GSR = "ENABLED";
    FD1P3IX timeout_count__i28 (.D(n657[28]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i28.GSR = "ENABLED";
    FD1P3IX timeout_count__i29 (.D(n657[29]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i29.GSR = "ENABLED";
    FD1P3IX timeout_count__i30 (.D(n657[30]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i30.GSR = "ENABLED";
    FD1P3IX timeout_count__i31 (.D(n657[31]), .SP(n9368), .CD(n9580), 
            .CK(debug_c_c), .Q(timeout_count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i31.GSR = "ENABLED";
    CCU2D add_30_11 (.A0(timeout_count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26423), .COUT(n26424), .S0(n657[9]), .S1(n657[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_11.INIT0 = 16'h5aaa;
    defparam add_30_11.INIT1 = 16'h5aaa;
    defparam add_30_11.INJECT1_0 = "NO";
    defparam add_30_11.INJECT1_1 = "NO";
    CCU2D add_30_27 (.A0(timeout_count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26431), .COUT(n26432), .S0(n657[25]), 
          .S1(n657[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_27.INIT0 = 16'h5aaa;
    defparam add_30_27.INIT1 = 16'h5aaa;
    defparam add_30_27.INJECT1_0 = "NO";
    defparam add_30_27.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_4_lut (.A(n31511), .B(register_addr[1]), .C(n31476), 
         .D(n31442), .Z(n29136)) /* synthesis lut_function=(A (B)+!A !((C (D))+!B)) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h8ccc;
    LUT4 i14485_3_lut (.A(Stepper_Y_Dir_c), .B(div_factor_reg_adj_993[5]), 
         .C(register_addr[1]), .Z(n21219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14485_3_lut.init = 16'hcaca;
    FD1P3AX reset_count_2668_2669__i2 (.D(n33690[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i2.GSR = "ENABLED";
    LUT4 i14477_3_lut (.A(Stepper_Y_En_c), .B(div_factor_reg_adj_993[6]), 
         .C(register_addr[1]), .Z(n21211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14477_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_281_4_lut_4_lut (.A(n31511), .B(n31476), .C(prev_select), 
         .D(n31473), .Z(n31424)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_rep_281_4_lut_4_lut.init = 16'h0400;
    LUT4 i14474_3_lut (.A(control_reg_adj_992[3]), .B(div_factor_reg_adj_993[3]), 
         .C(register_addr[1]), .Z(n21208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14474_3_lut.init = 16'hcaca;
    CCU2D add_30_25 (.A0(timeout_count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26430), .COUT(n26431), .S0(n657[23]), 
          .S1(n657[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_25.INIT0 = 16'h5aaa;
    defparam add_30_25.INIT1 = 16'h5aaa;
    defparam add_30_25.INJECT1_0 = "NO";
    defparam add_30_25.INJECT1_1 = "NO";
    CCU2D add_30_23 (.A0(timeout_count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26429), .COUT(n26430), .S0(n657[21]), 
          .S1(n657[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_23.INIT0 = 16'h5aaa;
    defparam add_30_23.INIT1 = 16'h5aaa;
    defparam add_30_23.INJECT1_0 = "NO";
    defparam add_30_23.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_511 (.A(n31511), .B(prev_select_adj_694), 
         .C(n31469), .D(select[4]), .Z(n14650)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_511.init = 16'h1000;
    FD1P3AX reset_count_2668_2669__i3 (.D(n33690[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i4 (.D(n33690[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i5 (.D(n33690[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i6 (.D(n33690[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i7 (.D(n33690[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i8 (.D(n33690[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i9 (.D(n33690[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i10 (.D(n33690[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i11 (.D(n33690[10]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i12 (.D(n33690[11]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i13 (.D(n33690[12]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i14 (.D(n33690[13]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2668_2669__i15 (.D(n33690[14]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669__i15.GSR = "ENABLED";
    CCU2D add_30_21 (.A0(timeout_count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26428), .COUT(n26429), .S0(n657[19]), 
          .S1(n657[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_21.INIT0 = 16'h5aaa;
    defparam add_30_21.INIT1 = 16'h5aaa;
    defparam add_30_21.INJECT1_0 = "NO";
    defparam add_30_21.INJECT1_1 = "NO";
    CCU2D reset_count_2668_2669_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n26889), .S0(n33690[13]), 
          .S1(n33690[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2668_2669_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n26888), .COUT(n26889), .S0(n33690[11]), 
          .S1(n33690[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2668_2669_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n26887), .COUT(n26888), .S0(n33690[9]), 
          .S1(n33690[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2668_2669_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n26886), .COUT(n26887), .S0(n33690[7]), 
          .S1(n33690[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_9.INJECT1_1 = "NO";
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.read_value({read_value_adj_1034}), 
            .debug_c_c(debug_c_c), .n2846(n2846), .GND_net(GND_net), .VCC_net(VCC_net), 
            .Stepper_Z_nFault_c(Stepper_Z_nFault_c), .n31511(n31511), .\read_size[0] (read_size_adj_1035[0]), 
            .n27752(n27752), .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n31419(n31419), 
            .databus({databus}), .limit_latched(limit_latched_adj_702), 
            .prev_limit_latched(prev_limit_latched_adj_703), .n9304(n9304), 
            .prev_select(prev_select_adj_738), .n31482(n31482), .\read_size[2] (read_size_adj_1035[2]), 
            .n29300(n29300), .\register_addr[1] (register_addr[1]), .\register_addr[5] (register_addr[5]), 
            .n31496(n31496), .rw(rw), .\select[4] (select[4]), .n52(n52_adj_695), 
            .\read_size[0]_adj_312 (read_size_adj_996[0]), .n5(n5), .prev_select_adj_313(prev_select_adj_694), 
            .n31421(n31421), .\steps_reg[7] (steps_reg_adj_1033[7]), .n31600(n31600), 
            .n31555(n31555), .n31590(n31590), .n31595(n31595), .\register_addr[4] (register_addr[4]), 
            .n29270(n29270), .n31463(n31463), .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), 
            .\register_addr[0] (register_addr[0]), .n29234(n29234), .n31503(n31503), 
            .\read_size[2]_adj_314 (read_size_adj_984[2]), .n9(n9_adj_899), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .n14522(n14522), .n610(n580_adj_1053[2]), 
            .n608(n580_adj_1053[4]), .Stepper_Z_Dir_c(Stepper_Z_Dir_c), 
            .Stepper_Z_En_c(Stepper_Z_En_c), .n11208(n11208), .n14546(n14546), 
            .\register_addr[3] (register_addr[3]), .\register_addr[2] (register_addr[2]), 
            .n31540(n31540), .n6(n33623[0]), .n4006(n4006), .Stepper_Z_Step_c(Stepper_Z_Step_c), 
            .limit_c_2(limit_c_2), .n11(n11), .n31410(n31410), .n16841(n16841), 
            .n8263(n8263), .n8297(n8297)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(608[25] 621[45])
    LUT4 i3_4_lut_4_lut (.A(n31511), .B(n31555), .C(n31595), .D(n29236), 
         .Z(n35)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_4_lut.init = 16'h0100;
    CCU2D reset_count_2668_2669_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n26885), .COUT(n26886), .S0(n33690[5]), 
          .S1(n33690[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_7.INJECT1_1 = "NO";
    CCU2D reset_count_2668_2669_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n26884), .COUT(n26885), .S0(n33690[3]), 
          .S1(n33690[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_5.INJECT1_1 = "NO";
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.debug_c_c(debug_c_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .n31511(n31511), .n4094({n4094}), .\read_size[0] (read_size_adj_996[0]), 
            .n14650(n14650), .n27751(n27751), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), 
            .databus({databus}), .prev_step_clk(prev_step_clk_adj_659), 
            .step_clk(step_clk_adj_658), .limit_latched(limit_latched_adj_656), 
            .prev_limit_latched(prev_limit_latched_adj_657), .n9300(n9300), 
            .prev_select(prev_select_adj_694), .n31445(n31445), .n29270(n29270), 
            .n29491(n29491), .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), .\register_addr[0] (register_addr[0]), 
            .\div_factor_reg[9] (div_factor_reg_adj_993[9]), .\div_factor_reg[6] (div_factor_reg_adj_993[6]), 
            .\div_factor_reg[5] (div_factor_reg_adj_993[5]), .\div_factor_reg[4] (div_factor_reg_adj_993[4]), 
            .\div_factor_reg[3] (div_factor_reg_adj_993[3]), .\control_reg[7] (control_reg_adj_992[7]), 
            .n12148(n12148), .Stepper_Y_En_c(Stepper_Y_En_c), .Stepper_Y_Dir_c(Stepper_Y_Dir_c), 
            .\control_reg[4] (control_reg_adj_992[4]), .\control_reg[3] (control_reg_adj_992[3]), 
            .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), .\read_size[2] (read_size_adj_996[2]), 
            .n29199(n29199), .\steps_reg[9] (steps_reg_adj_994[9]), .\steps_reg[6] (steps_reg_adj_994[6]), 
            .\steps_reg[5] (steps_reg_adj_994[5]), .\steps_reg[4] (steps_reg_adj_994[4]), 
            .\steps_reg[3] (steps_reg_adj_994[3]), .read_value({read_value_adj_995}), 
            .n9547(n9547), .\register_addr[1] (register_addr[1]), .n29112(n29112), 
            .limit_c_1(limit_c_1), .int_step(int_step), .n22(n22), .n31418(n31418), 
            .n29113(n29113), .n21213(n21213), .n21221(n21221), .n28826(n28826), 
            .n6807(n6778[3]), .n32(n32_adj_619), .n27483(n27483), .n224({n224_adj_999}), 
            .n8635(n8634[7]), .n8193(n8193), .n31407(n31407), .n16840(n16840), 
            .n8159(n8159)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(593[25] 606[45])
    CCU2D reset_count_2668_2669_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n26883), .COUT(n26884), .S0(n33690[1]), 
          .S1(n33690[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2668_2669_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2668_2669_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26883), .S1(n33690[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2668_2669_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2668_2669_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2668_2669_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2668_2669_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(register_addr[1]), .B(n9547), .Z(n29112)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut.init = 16'h2222;
    RCPeripheral rc_receiver (.n2(n2_adj_925), .databus({databus}), .\read_value[10] (read_value_adj_1073[10]), 
            .n8(n8_adj_927), .n31425(n31425), .\register_addr[0] (register_addr[0]), 
            .read_value({read_value}), .read_value_adj_308({read_value_adj_983}), 
            .n46(n46), .n52(n52), .databus_out({databus_out}), .rw(rw), 
            .read_value_adj_309({read_value_adj_995}), .\read_value[10]_adj_157 (read_value_adj_1119[10]), 
            .n52_adj_158(n52_adj_695), .n31446(n31446), .n2_adj_159(n2_adj_929), 
            .\read_value[9]_adj_160 (read_value_adj_1073[9]), .n8_adj_161(n8_adj_931), 
            .\read_value[9]_adj_162 (read_value_adj_1119[9]), .n2_adj_163(n2_adj_926), 
            .\select[7] (select[7]), .n176(n176), .\read_value[8]_adj_164 (read_value_adj_1073[8]), 
            .n8_adj_165(n8_adj_928), .\register_addr[1] (register_addr[1]), 
            .n2_adj_166(n2_adj_937), .\read_value[24]_adj_167 (read_value_adj_1073[24]), 
            .n8_adj_168(n8), .\read_value[24]_adj_169 (read_value_adj_1119[24]), 
            .\read_value[8]_adj_170 (read_value_adj_1119[8]), .n2_adj_171(n2_adj_930), 
            .\read_value[7]_adj_172 (read_value_adj_1119[7]), .\read_value[7]_adj_173 (read_value_adj_1111[7]), 
            .n31443(n31443), .n3(n3_adj_932), .read_value_adj_310({read_value_adj_976}), 
            .n64(n64), .n66(n66), .read_value_adj_311({read_value_adj_1135}), 
            .\read_value[14]_adj_190 (read_value_adj_1119[14]), .n2_adj_191(n2_adj_741), 
            .\read_value[6]_adj_192 (read_value_adj_1119[6]), .\read_value[6]_adj_193 (read_value_adj_1111[6]), 
            .n3_adj_194(n3_adj_948), .n2_adj_195(n2_adj_606), .\read_value[5]_adj_196 (read_value_adj_1119[5]), 
            .\read_value[5]_adj_197 (read_value_adj_1111[5]), .n33384(n33384), 
            .n3_adj_198(n3), .n2_adj_199(n2_adj_902), .\read_value[4]_adj_200 (read_value_adj_1119[4]), 
            .\read_value[4]_adj_201 (read_value_adj_1111[4]), .n3_adj_202(n3_adj_901), 
            .n2_adj_203(n2_adj_817), .\read_value[3]_adj_204 (read_value_adj_1119[3]), 
            .\read_value[3]_adj_205 (read_value_adj_1111[3]), .n2_adj_206(n2_adj_900), 
            .\read_value[22]_adj_207 (read_value_adj_1073[22]), .n8_adj_208(n8_adj_740), 
            .n3_adj_209(n3_adj_947), .n2_adj_210(n2_adj_936), .\read_value[2]_adj_211 (read_value_adj_1119[2]), 
            .\read_value[2]_adj_212 (read_value_adj_1111[2]), .\read_value[22]_adj_213 (read_value_adj_1119[22]), 
            .n3_adj_214(n3_adj_620), .n10(n10), .\read_value[1]_adj_215 (read_value_adj_1111[1]), 
            .n3_adj_216(n3_adj_701), .\read_value[1]_adj_217 (read_value_adj_1073[1]), 
            .n2_adj_218(n2_adj_923), .\read_value[13]_adj_219 (read_value_adj_1073[13]), 
            .n8_adj_220(n8_adj_924), .n2_adj_221(n2_adj_742), .\read_value[13]_adj_222 (read_value_adj_1119[13]), 
            .\read_value[23]_adj_223 (read_value_adj_1073[23]), .n8_adj_224(n8_adj_739), 
            .n2_adj_225(n2_adj_700), .n2_adj_226(n2_adj_933), .\read_value[12]_adj_227 (read_value_adj_1073[12]), 
            .n8_adj_228(n8_adj_935), .\read_value[23]_adj_229 (read_value_adj_1119[23]), 
            .\read_value[12]_adj_230 (read_value_adj_1119[12]), .\read_value[21]_adj_231 (read_value_adj_1073[21]), 
            .n8_adj_232(n8_adj_945), .read_size({read_size}), .\select[1] (select[1]), 
            .n13(n13_adj_699), .n31482(n31482), .n9(n9), .\read_size[0]_adj_233 (read_size_adj_1035[0]), 
            .n18(n18), .\read_size[0]_adj_234 (read_size_adj_1112[0]), .\read_size[0]_adj_235 (read_size_adj_977[0]), 
            .n31464(n31464), .\select[2] (select[2]), .n14(n14_adj_698), 
            .n31473(n31473), .n5(n5), .\read_size[0]_adj_236 (read_size_adj_984[0]), 
            .\read_size[0]_adj_237 (read_size_adj_1136[0]), .n31444(n31444), 
            .\select[5] (select[5]), .\read_size[0]_adj_238 (read_size_adj_1074[0]), 
            .n2_adj_239(n2), .\read_value[11]_adj_240 (read_value_adj_1073[11]), 
            .n8_adj_241(n8_adj_608), .n6(n6), .\read_size[2]_adj_242 (read_size_adj_1074[2]), 
            .\reg_size[2] (reg_size[2]), .\read_size[2]_adj_243 (read_size_adj_1035[2]), 
            .n9_adj_244(n9_adj_899), .\read_size[2]_adj_245 (read_size_adj_1120[2]), 
            .n31470(n31470), .\read_value[11]_adj_246 (read_value_adj_1119[11]), 
            .\read_value[21]_adj_247 (read_value_adj_1119[21]), .n2_adj_248(n2_adj_609), 
            .\read_value[25]_adj_249 (read_value_adj_1073[25]), .n8_adj_250(n8_adj_697), 
            .\read_value[25]_adj_251 (read_value_adj_1119[25]), .\register_addr[2] (register_addr[2]), 
            .n2_adj_252(n2_adj_942), .n2_adj_253(n2_adj_915), .\read_value[20]_adj_254 (read_value_adj_1073[20]), 
            .n8_adj_255(n8_adj_946), .\read_value[16]_adj_256 (read_value_adj_1073[16]), 
            .n8_adj_257(n8_adj_916), .n31587(n31587), .\sendcount[1] (sendcount[1]), 
            .n13155(n13155), .n31456(n31456), .\read_value[20]_adj_258 (read_value_adj_1119[20]), 
            .n2_adj_259(n2_adj_921), .n2_adj_260(n2_adj_605), .\read_value[0]_adj_261 (read_value_adj_1119[0]), 
            .\read_value[0]_adj_262 (read_value_adj_1111[0]), .n3_adj_263(n3_adj_607), 
            .n2_adj_264(n2_adj_914), .\read_value[26]_adj_265 (read_value_adj_1073[26]), 
            .n8_adj_266(n8_adj_913), .\read_value[26]_adj_267 (read_value_adj_1119[26]), 
            .\read_value[16]_adj_268 (read_value_adj_1119[16]), .n2_adj_269(n2_adj_943), 
            .\read_value[19]_adj_270 (read_value_adj_1073[19]), .n8_adj_271(n8_adj_818), 
            .n29236(n29236), .n2_adj_272(n2_adj_918), .\read_value[19]_adj_273 (read_value_adj_1119[19]), 
            .n2_adj_274(n2_adj_934), .\read_value[18]_adj_275 (read_value_adj_1073[18]), 
            .n8_adj_276(n8_adj_813), .n2_adj_277(n2_adj_903), .\read_value[31]_adj_278 (read_value_adj_1073[31]), 
            .n8_adj_279(n8_adj_904), .\read_value[14]_adj_280 (read_value_adj_1073[14]), 
            .n8_adj_281(n8_adj_922), .\read_value[31]_adj_282 (read_value_adj_1119[31]), 
            .n2_adj_283(n2_adj_816), .\read_value[30]_adj_284 (read_value_adj_1073[30]), 
            .n8_adj_285(n8_adj_906), .\read_value[18]_adj_286 (read_value_adj_1119[18]), 
            .\read_value[30]_adj_287 (read_value_adj_1119[30]), .n2_adj_288(n2_adj_908), 
            .\read_value[17]_adj_289 (read_value_adj_1119[17]), .\read_value[29]_adj_290 (read_value_adj_1073[29]), 
            .n8_adj_291(n8_adj_815), .\read_value[29]_adj_292 (read_value_adj_1119[29]), 
            .n2_adj_293(n2_adj_911), .n2_adj_294(n2_adj_917), .\read_value[15]_adj_295 (read_value_adj_1073[15]), 
            .n8_adj_296(n8_adj_920), .\read_value[28]_adj_297 (read_value_adj_1073[28]), 
            .n8_adj_298(n8_adj_909), .\read_value[17]_adj_299 (read_value_adj_1073[17]), 
            .n8_adj_300(n8_adj_919), .\read_value[28]_adj_301 (read_value_adj_1119[28]), 
            .n2_adj_302(n2_adj_912), .\read_value[27]_adj_303 (read_value_adj_1073[27]), 
            .n8_adj_304(n8_adj_814), .\read_value[15]_adj_305 (read_value_adj_1119[15]), 
            .\read_value[27]_adj_306 (read_value_adj_1119[27]), .GND_net(GND_net), 
            .debug_c_c(debug_c_c), .n33386(n33386), .rc_ch8_c(rc_ch8_c), 
            .n29817(n29817), .n33385(n33385), .n13956(n13956), .n27563(n27563), 
            .n29783(n29783), .rc_ch7_c(rc_ch7_c), .n33387(n33387), .n27542(n27542), 
            .n29826(n29826), .rc_ch4_c(rc_ch4_c), .n27549(n27549), .n29837(n29837), 
            .rc_ch3_c(rc_ch3_c), .n14499(n14499), .n27540(n27540), .n29839(n29839), 
            .n29529(n29529), .n29943(n29943), .n14_adj_307(n14_adj_910), 
            .n29831(n29831), .rc_ch2_c(rc_ch2_c), .n31411(n31411), .n14512(n14512), 
            .n29846(n29846), .n27535(n27535), .n31511(n31511), .n14513(n14513), 
            .rc_ch1_c(rc_ch1_c), .n29829(n29829), .n27546(n27546), .n29810(n29810)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(706[15] 718[41])
    LUT4 i15745_1_lut_rep_471 (.A(reset_count[14]), .B(reset_count[12]), 
         .C(reset_count[13]), .D(n29263), .Z(n33389)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam i15745_1_lut_rep_471.init = 16'h0515;
    SabertoothSerialPeripheral motor_serial (.\read_size[0] (read_size_adj_977[0]), 
            .debug_c_c(debug_c_c), .n9378(n9378), .n13907(n13907), .n31511(n31511), 
            .\databus[0] (databus[0]), .\select[2] (select[2]), .read_value({read_value_adj_976}), 
            .n9541(n9541), .rw(rw), .n64(n64), .n31600(n31600), .\register[0][7] (\register[0]_adj_975 [7]), 
            .n31581(n31581), .\reset_count[14] (reset_count[14]), .n22483(n22483), 
            .n11235(n11235), .\databus[7] (databus[7]), .\databus[6] (databus[6]), 
            .\databus[5] (databus[5]), .\databus[4] (databus[4]), .\databus[3] (databus[3]), 
            .\databus[2] (databus[2]), .\databus[1] (databus[1]), .\register_addr[0] (register_addr[0]), 
            .n31412(n31412), .GND_net(GND_net), .n1155(n1155), .n31536(n31536), 
            .\reset_count[8] (reset_count[8]), .\reset_count[7] (reset_count[7]), 
            .n29331(n29331), .state({state_adj_1312}), .n29169(n29169), 
            .n31595(n31595), .n31555(n31555), .n31575(n31575), .n9(n9_adj_938), 
            .n33384(n33384), .n31442(n31442), .n31589(n31589), .n35(n35), 
            .n4180(n4180), .\register_addr[5] (register_addr[5]), .n31463(n31463), 
            .n13916(n13916), .\reset_count[11] (reset_count[11]), .n21502(n21502), 
            .n27249(n27249), .n29263(n29263), .n14782(n14782), .n31529(n31529), 
            .n9296(n9296), .n31462(n31462), .motor_pwm_l_c(motor_pwm_l_c), 
            .n8506(n8506), .n29785(n29785), .select_clk(select_clk), .n2966(n2966), 
            .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(528[29] 536[56])
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 Select_4240_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[24]), 
         .D(rw), .Z(n8)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4240_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    \ProtocolInterface(baud_div=12)  protocol_interface (.register_addr({Open_0, 
            Open_1, register_addr[5:0]}), .debug_c_c(debug_c_c), .databus({databus}), 
            .\select[7] (select[7]), .n33389(n33389), .\select[5] (select[5]), 
            .\select[4] (select[4]), .\select[3] (select[3]), .\select[2] (select[2]), 
            .\select[1] (select[1]), .databus_out({databus_out}), .n13833(n13833), 
            .\sendcount[1] (sendcount[1]), .n31555(n31555), .n29300(n29300), 
            .n31532(n31532), .n29199(n29199), .debug_c_5(debug_c_5), .n31496(n31496), 
            .rw(rw), .n31425(n31425), .prev_select(prev_select_adj_780), 
            .n31427(n31427), .n31595(n31595), .n31469(n31469), .n31465(n31465), 
            .n31426(n31426), .\register[1][19] (\register[1]_adj_1109 [19]), 
            .n59(n99_adj_1336[19]), .n31500(n31500), .\register[1][20] (\register[1]_adj_1109 [20]), 
            .n57(n99_adj_1336[20]), .\register[1][26] (\register[1]_adj_1109 [26]), 
            .n45(n99_adj_1336[26]), .force_pause(force_pause), .\register[2] ({\register[2] }), 
            .\register[1][0] (\register[1]_adj_1109 [0]), .n97(n99_adj_1336[0]), 
            .n31503(n31503), .prev_select_adj_5(prev_select), .n31511(n31511), 
            .n13940(n13940), .n1491(n1473[14]), .n29169(n29169), .n29294(n29294), 
            .n29068(n29068), .n29292(n29292), .n31435(n31435), .n303(n303), 
            .n56(n56), .n29293(n29293), .n29065(n29065), .n29055(n29055), 
            .n29052(n29052), .n29064(n29064), .n29062(n29062), .n29049(n29049), 
            .n224({n224_adj_1077}), .n3921({n3921}), .n29051(n29051), 
            .n29053(n29053), .n27751(n27751), .n29066(n29066), .n29056(n29056), 
            .n29067(n29067), .n29070(n29070), .n29071(n29071), .n27752(n27752), 
            .n29069(n29069), .n29057(n29057), .n29058(n29058), .n29063(n29063), 
            .n29059(n29059), .n29257(n29257), .n29061(n29061), .n29054(n29054), 
            .n29050(n29050), .n29048(n29048), .n29060(n29060), .n29047(n29047), 
            .prev_select_adj_6(prev_select_adj_738), .n2846(n2846), .n66(n66), 
            .\register[0][2] (\register[0] [2]), .read_value({read_value_adj_1034}), 
            .n33384(n33384), .n2(n2_adj_742), .n31464(n31464), .n2_adj_7(n2_adj_900), 
            .n2_adj_8(n2_adj_700), .n2_adj_9(n2_adj_942), .n2_adj_10(n2_adj_609), 
            .n31540(n31540), .n31449(n31449), .n31477(n31477), .n31470(n31470), 
            .n2_adj_11(n2_adj_937), .n2_adj_12(n2_adj_943), .n2_adj_13(n2_adj_934), 
            .n31473(n31473), .n2_adj_14(n2_adj_917), .n2_adj_15(n2_adj_915), 
            .n2_adj_16(n2_adj_918), .n2_adj_17(n2_adj_921), .n2_adj_18(n2_adj_923), 
            .n2_adj_19(n2_adj_933), .n2_adj_20(n2), .n2_adj_21(n2_adj_925), 
            .n2_adj_22(n2_adj_929), .n2_adj_23(n2_adj_926), .n3(n3_adj_932), 
            .n3_adj_24(n3_adj_948), .n3_adj_25(n3), .n31589(n31589), .n31476(n31476), 
            .n3_adj_26(n3_adj_901), .n3_adj_27(n3_adj_947), .n3_adj_28(n3_adj_620), 
            .n3_adj_29(n3_adj_701), .n3_adj_30(n3_adj_607), .n2_adj_31(n2_adj_903), 
            .n2_adj_32(n2_adj_816), .n2_adj_33(n2_adj_908), .n2_adj_34(n2_adj_911), 
            .n2_adj_35(n2_adj_912), .n2_adj_36(n2_adj_914), .n31482(n31482), 
            .n14453(n14453), .n9537(n9537), .n35(n35), .n27464(n27464), 
            .n33383(n33383), .n31445(n31445), .debug_c_7(debug_c_7), .\read_size[2] (read_size_adj_996[2]), 
            .n29234(n29234), .n31444(n31444), .n52(n52), .n31442(n31442), 
            .n29236(n29236), .n176(n176), .n31448(n31448), .n31570(n31570), 
            .n16012(n16012), .n31456(n31456), .n31581(n31581), .n13907(n13907), 
            .n11235(n11235), .n31434(n31434), .n30305(n30305), .n29220(n29220), 
            .n31525(n31525), .n31419(n31419), .n30303(n30303), .\control_reg[7] (control_reg[7]), 
            .n1(n1), .n31529(n31529), .n31539(n31539), .n13155(n13155), 
            .n13(n13_adj_699), .n18(n18), .n14(n14_adj_698), .\reg_size[2] (reg_size[2]), 
            .n31587(n31587), .n31590(n31590), .n27441(n27441), .\control_reg[7]_adj_37 (control_reg_adj_1070[7]), 
            .n31600(n31600), .n32(n32), .n4(n4), .n5833(n5833), .prev_select_adj_38(prev_select_adj_898), 
            .\reset_count[14] (reset_count[14]), .n22483(n22483), .n2869(n2869), 
            .n224_adj_91({n224_adj_999}), .n4094({n4094}), .n31575(n31575), 
            .\read_value[7]_adj_71 (read_value_adj_1073[7]), .n2_adj_72(n2_adj_930), 
            .\read_value[5]_adj_73 (read_value_adj_1073[5]), .n2_adj_74(n2_adj_606), 
            .n31472(n31472), .\read_value[4]_adj_75 (read_value_adj_1073[4]), 
            .n2_adj_76(n2_adj_902), .\read_value[6]_adj_77 (read_value_adj_1073[6]), 
            .n2_adj_78(n2_adj_741), .\read_value[3]_adj_79 (read_value_adj_1073[3]), 
            .n2_adj_80(n2_adj_817), .\read_value[2]_adj_81 (read_value_adj_1073[2]), 
            .n2_adj_82(n2_adj_936), .\read_value[0]_adj_83 (read_value_adj_1073[0]), 
            .n2_adj_84(n2_adj_605), .n27444(n27444), .n34(n34), .n29256(n29256), 
            .n9330(n9330), .n1485(n1473[20]), .\register[0][5] (\register[0]_adj_1134 [5]), 
            .expansion5_c(expansion5_c), .\register[1][5] (\register[1]_adj_1133 [5]), 
            .debug_c_2(debug_c_2), .n1488(n1473[17]), .debug_c_3(debug_c_3), 
            .n9378(n9378), .n29491(n29491), .prev_select_adj_85(prev_select_adj_694), 
            .\steps_reg[7] (steps_reg_adj_1033[7]), .n11(n11), .debug_c_4(debug_c_4), 
            .n31501(n31501), .n6005(n5973[0]), .\steps_reg[5] (steps_reg_adj_994[5]), 
            .n14_adj_86(n14), .\register[0][4] (\register[0]_adj_1134 [4]), 
            .expansion4_out(expansion4_out), .\register[1][4] (\register[1]_adj_1133 [4]), 
            .timeout_pause(timeout_pause), .\steps_reg[6] (steps_reg_adj_994[6]), 
            .n13_adj_87(n13), .\register[0][7] (\register[0]_adj_975 [7]), 
            .n31536(n31536), .clk_1Hz(clk_1Hz), .signal_light_c(signal_light_c), 
            .\steps_reg[3] (steps_reg_adj_994[3]), .n12(n12), .\control_reg[4] (control_reg_adj_992[4]), 
            .\div_factor_reg[4] (div_factor_reg_adj_993[4]), .\steps_reg[4] (steps_reg_adj_994[4]), 
            .\control_reg[7]_adj_88 (control_reg_adj_992[7]), .n8635(n8634[7]), 
            .n13947(n13947), .n12368(n12368), .n9300(n9300), .n14522(n14522), 
            .n4006(n4006), .n31406(n31406), .n27679(n27679), .n27483(n27483), 
            .n32_adj_89(n32_adj_619), .n16764(n16764), .n9(n9_adj_938), 
            .n9304(n9304), .prev_select_adj_90(prev_select_adj_853), .n16763(n16763), 
            .n6002(n5973[3]), .n27427(n27427), .n28826(n28826), .n8653(n8652[7]), 
            .\state[3] (state_adj_1312[3]), .\state[1] (state_adj_1312[1]), 
            .\state[0] (state_adj_1312[0]), .n1155(n1155), .n73(n73), 
            .\reset_count[7] (reset_count[7]), .\reset_count[6] (reset_count[6]), 
            .\reset_count[5] (reset_count[5]), .n27249(n27249), .n11072(n11072), 
            .GND_net(GND_net), .uart_rx_c(uart_rx_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(493[26] 503[57])
    CCU2D add_30_19 (.A0(timeout_count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26427), .COUT(n26428), .S0(n657[17]), 
          .S1(n657[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_30_19.INIT0 = 16'h5aaa;
    defparam add_30_19.INIT1 = 16'h5aaa;
    defparam add_30_19.INJECT1_0 = "NO";
    defparam add_30_19.INJECT1_1 = "NO";
    LUT4 Select_4237_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[25]), 
         .D(rw), .Z(n8_adj_697)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4237_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4243_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[23]), 
         .D(rw), .Z(n8_adj_739)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4243_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4246_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[22]), 
         .D(rw), .Z(n8_adj_740)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4246_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4249_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[21]), 
         .D(rw), .Z(n8_adj_945)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4249_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2657_1_lut (.A(n7846), .Z(n9368)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2657_1_lut.init = 16'h5555;
    LUT4 i29_2_lut (.A(uart_rx_c), .B(prev_uart_rx), .Z(n9580)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[7:29])
    defparam i29_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_512 (.A(div_factor_reg_adj_993[9]), .B(n29112), .C(steps_reg_adj_994[9]), 
         .D(register_addr[0]), .Z(n29113)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_512.init = 16'hc088;
    LUT4 Select_4252_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[20]), 
         .D(rw), .Z(n8_adj_946)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4252_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4255_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[19]), 
         .D(rw), .Z(n8_adj_818)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4255_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i14487 (.BLUT(n21219), .ALUT(n14), .C0(register_addr[0]), .Z(n21221));
    LUT4 Select_4258_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[18]), 
         .D(rw), .Z(n8_adj_813)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4258_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4261_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[17]), 
         .D(rw), .Z(n8_adj_919)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4261_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4264_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[16]), 
         .D(rw), .Z(n8_adj_916)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4264_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i22314_2_lut (.A(int_step), .B(control_reg_adj_992[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i22314_2_lut.init = 16'h9999;
    LUT4 Select_4267_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[15]), 
         .D(rw), .Z(n8_adj_920)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4267_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i14479 (.BLUT(n21211), .ALUT(n13), .C0(register_addr[0]), .Z(n21213));
    LUT4 Select_4270_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[14]), 
         .D(n33384), .Z(n8_adj_922)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4270_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    GlobalControlPeripheral global_control (.\register[2] ({\register[2] }), 
            .GND_net(GND_net), .force_pause(force_pause), .debug_c_c(debug_c_c), 
            .n31511(n31511), .\databus[1] (databus[1]), .n9483(n9483), 
            .read_size({read_size}), .n14453(n14453), .n31449(n31449), 
            .prev_clk_1Hz(prev_clk_1Hz), .clk_1Hz(clk_1Hz), .\register[0][2] (\register[0] [2]), 
            .\select[1] (select[1]), .read_value({read_value}), .n29068(n29068), 
            .rw(rw), .n46(n46), .n29292(n29292), .n31477(n31477), .n29293(n29293), 
            .n29294(n29294), .n30305(n30305), .n30303(n30303), .\reset_count[14] (reset_count[14]), 
            .n22483(n22483), .xbee_pause_c(xbee_pause_c), .\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .n29169(n29169), .n9537(n9537), 
            .n6002(n5973[3]), .n29065(n29065), .n29055(n29055), .n29052(n29052), 
            .n16764(n16764), .n27427(n27427), .n29064(n29064), .n16763(n16763), 
            .n29062(n29062), .n29049(n29049), .n29051(n29051), .n29053(n29053), 
            .n29066(n29066), .n29056(n29056), .n29067(n29067), .n29070(n29070), 
            .n29071(n29071), .n29069(n29069), .n6005(n5973[0]), .n29057(n29057), 
            .n29058(n29058), .n29063(n29063), .n29059(n29059), .n29061(n29061), 
            .n29054(n29054), .n29050(n29050), .n29048(n29048), .n29060(n29060), 
            .n29047(n29047), .n29788(n29788), .n2875(n2875)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(514[45] 525[74])
    ClockDivider_U10 pwm_clk_div (.clk_255kHz(clk_255kHz), .debug_c_c(debug_c_c), 
            .n241(n241), .GND_net(GND_net), .n7916(n7916), .n31511(n31511), 
            .n7881(n7881), .n29831(n29831), .n14512(n14512), .n29829(n29829), 
            .n14513(n14513), .n2823(n2823), .n29839(n29839), .n27540(n27540), 
            .n29846(n29846), .n27535(n27535), .n29817(n29817), .n13956(n13956), 
            .n29529(n29529), .n14(n14_adj_910), .n29943(n29943), .n14499(n14499), 
            .n29783(n29783), .n27563(n27563), .n29810(n29810), .n27546(n27546), 
            .n29826(n29826), .n27542(n27542), .n29837(n29837), .n27549(n27549)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(538[15] 541[41])
    LUT4 Select_4273_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[13]), 
         .D(rw), .Z(n8_adj_924)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4273_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i14476 (.BLUT(n21208), .ALUT(n12), .C0(register_addr[0]), .Z(n6778[3]));
    LUT4 Select_4276_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[12]), 
         .D(rw), .Z(n8_adj_935)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4276_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4279_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[11]), 
         .D(rw), .Z(n8_adj_608)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4279_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.debug_c_c(debug_c_c), .n31511(n31511), 
            .databus({databus}), .n4180(n4180), .\read_size[0] (read_size_adj_984[0]), 
            .n13940(n13940), .n9378(n9378), .Stepper_X_M0_c_0(Stepper_X_M0_c_0), 
            .n13916(n13916), .prev_step_clk(prev_step_clk), .step_clk(step_clk), 
            .limit_latched(limit_latched), .prev_limit_latched(prev_limit_latched), 
            .n9296(n9296), .prev_select(prev_select), .n31473(n31473), 
            .\register_addr[1] (register_addr[1]), .Stepper_X_Dir_c(Stepper_X_Dir_c), 
            .\register_addr[0] (register_addr[0]), .n1(n1), .Stepper_X_En_c(Stepper_X_En_c), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\control_reg[7] (control_reg[7]), 
            .n12158(n12158), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), .\read_size[2] (read_size_adj_984[2]), 
            .n31434(n31434), .n34(n34), .n27444(n27444), .n29136(n29136), 
            .limit_c_0(limit_c_0), .read_value({read_value_adj_983}), .n31424(n31424), 
            .n24(n24), .n31420(n31420), .VCC_net(VCC_net), .GND_net(GND_net), 
            .Stepper_X_nFault_c(Stepper_X_nFault_c), .Stepper_X_Step_c(Stepper_X_Step_c), 
            .n31408(n31408), .n8055(n8055), .n8089(n8089), .n17034(n17034)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(578[25] 591[45])
    LUT4 Select_4282_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[10]), 
         .D(n33384), .Z(n8_adj_927)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4282_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_4_lut (.A(n31511), .B(n303), .C(n31448), .D(n31570), 
         .Z(n24145)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h5400;
    LUT4 Select_4285_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[9]), 
         .D(n33384), .Z(n8_adj_931)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4285_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_4_lut_adj_513 (.A(n31511), .B(n31532), .C(n31539), .D(n31421), 
         .Z(n9547)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C+!(D))))) */ ;
    defparam i2_4_lut_4_lut_adj_513.init = 16'h4500;
    LUT4 Select_4288_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[8]), 
         .D(n33384), .Z(n8_adj_928)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4288_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4219_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[31]), 
         .D(n33384), .Z(n8_adj_904)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4219_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    EncoderPeripheral right_encoder (.\register_addr[0] (register_addr[0]), 
            .n31431(n31431), .prev_select(prev_select_adj_888), .debug_c_c(debug_c_c), 
            .n31470(n31470), .\read_size[0] (read_size_adj_1120[0]), .n15086(n15086), 
            .n6(n33623[0]), .encoder_rb_c(encoder_rb_c), .encoder_ra_c(encoder_ra_c), 
            .read_value({read_value_adj_1119}), .\read_size[2] (read_size_adj_1120[2]), 
            .n31540(n31540), .encoder_ri_c(encoder_ri_c), .qreset(qreset), 
            .VCC_net(VCC_net), .GND_net(GND_net), .\quadA_delayed[1] (quadA_delayed_adj_1223[1]), 
            .n13938(n13938), .n6_adj_4(n6_adj_944), .\quadB_delayed[1] (quadB_delayed_adj_1224[1])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(680[20] 690[47])
    \ClockDividerP_SP(factor=120000)  clk_100Hz_divider (.n29791(n29791), 
            .debug_c_0(debug_c_0), .debug_c_c(debug_c_c), .n31511(n31511), 
            .n2860(n2860), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(641[29] 643[61])
    LUT4 Select_4222_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[30]), 
         .D(n33384), .Z(n8_adj_906)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4222_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 m1_lut (.Z(n33383)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    LUT4 i15735_4_lut (.A(n22389), .B(n13315), .C(n21502), .D(n29331), 
         .Z(n22483)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i15735_4_lut.init = 16'hfcec;
    LUT4 i15646_3_lut (.A(reset_count[5]), .B(reset_count[6]), .C(reset_count[4]), 
         .Z(n22389)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15646_3_lut.init = 16'hc8c8;
    LUT4 Select_4225_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[29]), 
         .D(n33384), .Z(n8_adj_815)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4225_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    EncoderPeripheral_U11 left_encoder (.\read_size[0] (read_size_adj_1112[0]), 
            .debug_c_c(debug_c_c), .n14145(n14145), .n31426(n31426), .n31449(n31449), 
            .prev_select(prev_select_adj_853), .n31464(n31464), .\read_size[2] (read_size_adj_1112[2]), 
            .n31477(n31477), .read_value({read_value_adj_1111}), .\register_addr[0] (register_addr[0]), 
            .encoder_la_c(encoder_la_c), .encoder_lb_c(encoder_lb_c), .n59(n99_adj_1336[19]), 
            .n57(n99_adj_1336[20]), .n45(n99_adj_1336[26]), .\quadA_delayed[1] (quadA_delayed_adj_1223[1]), 
            .qreset(qreset), .n6(n6_adj_944), .\quadB_delayed[1] (quadB_delayed_adj_1224[1]), 
            .n13938(n13938), .n97(n99_adj_1336[0]), .encoder_li_c(encoder_li_c), 
            .GND_net(GND_net), .\register[1][0] (\register[1]_adj_1109 [0]), 
            .VCC_net(VCC_net), .\register[1][19] (\register[1]_adj_1109 [19]), 
            .\register[1][20] (\register[1]_adj_1109 [20]), .\register[1][26] (\register[1]_adj_1109 [26])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(669[20] 679[47])
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.read_value({read_value_adj_1073}), 
            .debug_c_c(debug_c_c), .n2857(n2857), .n31511(n31511), .n3921({n3921}), 
            .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_1074[0]), .n29257(n29257), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .databus({databus}), .limit_latched(limit_latched_adj_744), 
            .prev_limit_latched(prev_limit_latched_adj_745), .n9330(n9330), 
            .prev_select(prev_select_adj_780), .n31444(n31444), .Stepper_A_M1_c_1(Stepper_A_M1_c_1), 
            .\register_addr[0] (register_addr[0]), .\register_addr[1] (register_addr[1]), 
            .n224({n224_adj_1077}), .n32(n32), .n32_adj_1(n32_adj_619), 
            .prev_step_clk(prev_step_clk_adj_659), .step_clk(step_clk_adj_658), 
            .n31418(n31418), .n22(n22), .prev_step_clk_adj_2(prev_step_clk), 
            .n34(n34), .step_clk_adj_3(step_clk), .n31420(n31420), .n24(n24), 
            .n31427(n31427), .\register_addr[5] (register_addr[5]), .n31496(n31496), 
            .n29270(n29270), .n31575(n31575), .n27441(n27441), .\read_size[2] (read_size_adj_1074[2]), 
            .n29256(n29256), .Stepper_A_M2_c_2(Stepper_A_M2_c_2), .Stepper_A_Dir_c(Stepper_A_Dir_c), 
            .Stepper_A_En_c(Stepper_A_En_c), .\control_reg[7] (control_reg_adj_1070[7]), 
            .n12210(n12210), .Stepper_A_Step_c(Stepper_A_Step_c), .limit_c_3(limit_c_3), 
            .n8653(n8652[7]), .n31409(n31409), .n8401(n8401), .n8367(n8367), 
            .n16842(n16842)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(623[25] 636[45])
    LUT4 Select_4228_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31501), .C(read_value_adj_1111[28]), 
         .D(n33384), .Z(n8_adj_909)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(651[4] 667[11])
    defparam Select_4228_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    
endmodule
//
// Verilog Description of module ExpansionGPIO
//

module ExpansionGPIO (read_value, debug_c_c, n2869, n29220, n13947, 
            n31511, \databus[0] , \read_size[0] , n27679, prev_select, 
            \select[5] , expansion1_c_9, n31435, n56, expansion2_c_10, 
            expansion3_c_11, \databus[1] , \databus[2] , \databus[3] , 
            \register[0][4] , \databus[4] , \register[0][5] , \databus[5] , 
            \databus[6] , \databus[7] , n16012, \register[1][4] , \register[1][5] , 
            n12368, n31406, \register_addr[0] , n24145, n11007, n11006) /* synthesis syn_module_defined=1 */ ;
    output [7:0]read_value;
    input debug_c_c;
    input n2869;
    input n29220;
    input n13947;
    input n31511;
    input \databus[0] ;
    output \read_size[0] ;
    input n27679;
    output prev_select;
    input \select[5] ;
    output expansion1_c_9;
    input n31435;
    input n56;
    output expansion2_c_10;
    output expansion3_c_11;
    input \databus[1] ;
    input \databus[2] ;
    input \databus[3] ;
    output \register[0][4] ;
    input \databus[4] ;
    output \register[0][5] ;
    input \databus[5] ;
    input \databus[6] ;
    input \databus[7] ;
    input n16012;
    output \register[1][4] ;
    output \register[1][5] ;
    input n12368;
    input n31406;
    input \register_addr[0] ;
    input n24145;
    output n11007;
    output n11006;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]n7636;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]n7661;
    
    FD1P3AX read_value_i0_i4 (.D(n29220), .SP(n2869), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i4.GSR = "ENABLED";
    FD1P3IX register_0___i1 (.D(\databus[0] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i1.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n27679), .SP(n2869), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3AX prev_select_145 (.D(\select[5] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam prev_select_145.GSR = "ENABLED";
    LUT4 mux_2027_i2_4_lut (.A(expansion1_c_9), .B(\register[0] [1]), .C(n31435), 
         .D(n56), .Z(n7636[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2027_i2_4_lut.init = 16'ha0ac;
    LUT4 mux_2027_i3_4_lut (.A(expansion2_c_10), .B(\register[0] [2]), .C(n31435), 
         .D(n56), .Z(n7636[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2027_i3_4_lut.init = 16'ha0ac;
    LUT4 mux_2027_i4_4_lut (.A(expansion3_c_11), .B(\register[0] [3]), .C(n31435), 
         .D(n56), .Z(n7636[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2027_i4_4_lut.init = 16'ha0ac;
    FD1P3IX register_0___i2 (.D(\databus[1] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i2.GSR = "ENABLED";
    FD1P3IX register_0___i3 (.D(\databus[2] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i3.GSR = "ENABLED";
    FD1P3IX register_0___i4 (.D(\databus[3] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i4.GSR = "ENABLED";
    FD1P3IX register_0___i5 (.D(\databus[4] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i5.GSR = "ENABLED";
    FD1P3IX register_0___i6 (.D(\databus[5] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0][5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i6.GSR = "ENABLED";
    FD1P3IX register_0___i7 (.D(\databus[6] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i7.GSR = "ENABLED";
    FD1P3IX register_0___i8 (.D(\databus[7] ), .SP(n13947), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i8.GSR = "ENABLED";
    FD1P3IX register_0___i9 (.D(\databus[0] ), .SP(n16012), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i9.GSR = "ENABLED";
    FD1P3IX register_0___i10 (.D(\databus[1] ), .SP(n16012), .CD(n31511), 
            .CK(debug_c_c), .Q(expansion1_c_9)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i10.GSR = "ENABLED";
    FD1P3IX register_0___i11 (.D(\databus[2] ), .SP(n16012), .CD(n31511), 
            .CK(debug_c_c), .Q(expansion2_c_10)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i11.GSR = "ENABLED";
    FD1P3IX register_0___i12 (.D(\databus[3] ), .SP(n16012), .CD(n31511), 
            .CK(debug_c_c), .Q(expansion3_c_11)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i12.GSR = "ENABLED";
    FD1P3IX register_0___i13 (.D(\databus[4] ), .SP(n16012), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[1][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i13.GSR = "ENABLED";
    FD1P3IX register_0___i14 (.D(\databus[5] ), .SP(n16012), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[1][5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i14.GSR = "ENABLED";
    FD1P3IX register_0___i15 (.D(\databus[6] ), .SP(n16012), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i15.GSR = "ENABLED";
    FD1P3IX register_0___i16 (.D(\databus[7] ), .SP(n12368), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i16.GSR = "ENABLED";
    FD1P3AX read_value_i0_i1 (.D(n7636[1]), .SP(n2869), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i1.GSR = "ENABLED";
    FD1P3AX read_value_i0_i2 (.D(n7636[2]), .SP(n2869), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i2.GSR = "ENABLED";
    FD1P3AX read_value_i0_i3 (.D(n7636[3]), .SP(n2869), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i3.GSR = "ENABLED";
    FD1P3AX read_value_i0_i5 (.D(n31406), .SP(n2869), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i5.GSR = "ENABLED";
    LUT4 mux_2028_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n7661[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2028_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2028_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n7661[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2028_Mux_6_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value_i0_i7 (.D(n7661[7]), .SP(n2869), .CD(n24145), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i7.GSR = "ENABLED";
    FD1P3IX read_value_i0_i6 (.D(n7661[6]), .SP(n2869), .CD(n24145), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i6.GSR = "ENABLED";
    FD1P3IX read_value_i0_i0 (.D(n7661[0]), .SP(n2869), .CD(n24145), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=692, LSE_RLINE=703 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i0.GSR = "ENABLED";
    LUT4 mux_2028_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n7661[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2028_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 Select_4214_i3_4_lut (.A(\register[1][4] ), .B(\register[0][5] ), 
         .C(\register[0][4] ), .D(\register[1][5] ), .Z(n11007)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam Select_4214_i3_4_lut.init = 16'heca0;
    LUT4 i22468_2_lut (.A(\register[0][5] ), .B(\register[0][4] ), .Z(n11006)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22468_2_lut.init = 16'h1111;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (read_value, debug_c_c, n2846, 
            GND_net, VCC_net, Stepper_Z_nFault_c, n31511, \read_size[0] , 
            n27752, Stepper_Z_M0_c_0, n31419, databus, limit_latched, 
            prev_limit_latched, n9304, prev_select, n31482, \read_size[2] , 
            n29300, \register_addr[1] , \register_addr[5] , n31496, 
            rw, \select[4] , n52, \read_size[0]_adj_312 , n5, prev_select_adj_313, 
            n31421, \steps_reg[7] , n31600, n31555, n31590, n31595, 
            \register_addr[4] , n29270, n31463, Stepper_Z_M1_c_1, \register_addr[0] , 
            n29234, n31503, \read_size[2]_adj_314 , n9, Stepper_Z_M2_c_2, 
            n14522, n610, n608, Stepper_Z_Dir_c, Stepper_Z_En_c, n11208, 
            n14546, \register_addr[3] , \register_addr[2] , n31540, 
            n6, n4006, Stepper_Z_Step_c, limit_c_2, n11, n31410, 
            n16841, n8263, n8297) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2846;
    input GND_net;
    input VCC_net;
    input Stepper_Z_nFault_c;
    input n31511;
    output \read_size[0] ;
    input n27752;
    output Stepper_Z_M0_c_0;
    input n31419;
    input [31:0]databus;
    output limit_latched;
    output prev_limit_latched;
    input n9304;
    output prev_select;
    input n31482;
    output \read_size[2] ;
    input n29300;
    input \register_addr[1] ;
    input \register_addr[5] ;
    input n31496;
    input rw;
    input \select[4] ;
    output n52;
    input \read_size[0]_adj_312 ;
    output n5;
    input prev_select_adj_313;
    output n31421;
    output \steps_reg[7] ;
    input n31600;
    input n31555;
    output n31590;
    input n31595;
    input \register_addr[4] ;
    output n29270;
    output n31463;
    output Stepper_Z_M1_c_1;
    input \register_addr[0] ;
    input n29234;
    input n31503;
    input \read_size[2]_adj_314 ;
    output n9;
    output Stepper_Z_M2_c_2;
    input n14522;
    input n610;
    input n608;
    output Stepper_Z_Dir_c;
    output Stepper_Z_En_c;
    input n11208;
    input n14546;
    input \register_addr[3] ;
    input \register_addr[2] ;
    output n31540;
    output n6;
    input n4006;
    output Stepper_Z_Step_c;
    input limit_c_2;
    input n11;
    input n31410;
    input n16841;
    output n8263;
    output n8297;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n31616, n26845;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n224;
    
    wire n26846, n26844, n26843, n26842, fault_latched;
    wire [31:0]n4007;
    
    wire prev_step_clk, step_clk, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n31615, n31614, n26841, n26840, n26839, n26838, n26837, 
        n26836, n26835, n19910;
    wire [31:0]n100;
    
    wire n21, n17, n19, n19930, n29769, n29718, n27421;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n49, n62_adj_595, n58_adj_596, n50, n41, n60_adj_597, n54_adj_598, 
        n42_adj_599, n52_adj_600, n38_adj_601, n56_adj_602, n46_adj_603, 
        n29716, n29717, n27420, n29767, n29768, n19928;
    wire [7:0]n8643;
    
    wire int_step;
    wire [31:0]n7056;
    
    wire n10, n31417, n26850, n26849, n26848, n26847;
    
    FD1P3AX read_value__i0 (.D(n31616), .SP(n2846), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26845), .COUT(n26846), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26844), .COUT(n26845), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26843), .COUT(n26844), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26842), .COUT(n26843), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4007[0]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n27752), .SP(n2846), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n31419), .CD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31482), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n29300), .SP(n2846), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n4007[31]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4007[30]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4007[29]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4007[28]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4007[27]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4007[26]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4007[25]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    LUT4 n30929_bdd_4_lut_then_3_lut (.A(steps_reg[0]), .B(limit_latched), 
         .C(\register_addr[1] ), .Z(n31615)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n30929_bdd_4_lut_then_3_lut.init = 16'hacac;
    LUT4 n30929_bdd_4_lut_else_3_lut (.A(Stepper_Z_M0_c_0), .B(div_factor_reg[0]), 
         .C(\register_addr[1] ), .Z(n31614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30929_bdd_4_lut_else_3_lut.init = 16'hcaca;
    LUT4 i20_2_lut_3_lut_4_lut (.A(\register_addr[5] ), .B(n31496), .C(rw), 
         .D(\select[4] ), .Z(n52)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i20_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\register_addr[5] ), .B(n31496), .C(\read_size[0]_adj_312 ), 
         .D(\select[4] ), .Z(n5)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_278_3_lut_4_lut (.A(\register_addr[5] ), .B(n31496), 
         .C(prev_select_adj_313), .D(\select[4] ), .Z(n31421)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_278_3_lut_4_lut.init = 16'h0400;
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26841), .COUT(n26842), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26840), .COUT(n26841), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26839), .COUT(n26840), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(\steps_reg[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26838), .COUT(n26839), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26837), .COUT(n26838), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26836), .COUT(n26837), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26835), .COUT(n26836), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n19910), .D1(prev_step_clk), 
          .COUT(n26835), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n21), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n17), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n19), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n19930), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29769), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29718), .SP(n2846), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i2_3_lut (.A(n27421), .B(n31600), .C(control_reg[7]), .Z(n19910)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_3_lut.init = 16'h2020;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_595), .C(n58_adj_596), .D(n50), 
         .Z(n27421)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[15]), .B(steps_reg[23]), .C(steps_reg[21]), 
         .D(steps_reg[31]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_597), .C(n54_adj_598), .D(n42_adj_599), 
         .Z(n62_adj_595)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_504 (.A(n31555), .B(n31590), .C(n31595), 
         .D(\register_addr[4] ), .Z(n29270)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut_3_lut_4_lut_adj_504.init = 16'h0100;
    LUT4 i1_2_lut_rep_320_3_lut_4_lut (.A(n31555), .B(n31590), .C(n31595), 
         .D(\register_addr[4] ), .Z(n31463)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut_rep_320_3_lut_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[27]), .B(n52_adj_600), .C(n38_adj_601), 
         .D(steps_reg[20]), .Z(n58_adj_596)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[29]), .B(steps_reg[14]), .C(steps_reg[30]), 
         .D(steps_reg[19]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[16]), .B(steps_reg[24]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[8]), .B(n56_adj_602), .C(n46_adj_603), 
         .D(steps_reg[0]), .Z(n60_adj_597)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[9]), .B(steps_reg[17]), .C(steps_reg[12]), 
         .D(steps_reg[2]), .Z(n54_adj_598)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[25]), .B(steps_reg[26]), .Z(n42_adj_599)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[6]), .B(steps_reg[4]), .C(steps_reg[10]), 
         .D(steps_reg[3]), .Z(n56_adj_602)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[22]), .B(steps_reg[5]), .Z(n46_adj_603)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[13]), .B(steps_reg[18]), .C(steps_reg[28]), 
         .D(steps_reg[1]), .Z(n52_adj_600)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[11]), .B(\steps_reg[7] ), .Z(n38_adj_601)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i22156_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22156_3_lut.init = 16'hcaca;
    LUT4 i22157_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22157_3_lut.init = 16'hcaca;
    LUT4 i14896_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14896_4_lut.init = 16'hc088;
    LUT4 i14897_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14897_4_lut.init = 16'hc088;
    LUT4 i14898_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14898_4_lut.init = 16'hc088;
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[27]), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i14899_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14899_4_lut.init = 16'hc088;
    LUT4 i14900_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14900_4_lut.init = 16'hc088;
    LUT4 i14901_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14901_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_505 (.A(\register_addr[1] ), .B(div_factor_reg[23]), 
         .C(steps_reg[23]), .D(\register_addr[0] ), .Z(n21)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_505.init = 16'ha088;
    LUT4 i14902_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14902_4_lut.init = 16'hc088;
    LUT4 i14903_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14903_4_lut.init = 16'hc088;
    LUT4 i14904_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14904_4_lut.init = 16'hc088;
    LUT4 i14905_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14905_4_lut.init = 16'hc088;
    LUT4 i14906_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14906_4_lut.init = 16'hc088;
    LUT4 i14907_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14907_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_506 (.A(\register_addr[1] ), .B(div_factor_reg[16]), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n17)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_506.init = 16'ha088;
    LUT4 i1_4_lut_adj_507 (.A(\register_addr[1] ), .B(div_factor_reg[15]), 
         .C(steps_reg[15]), .D(\register_addr[0] ), .Z(n19)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_507.init = 16'ha088;
    LUT4 i14908_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14908_4_lut.init = 16'hc088;
    LUT4 i14909_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14909_4_lut.init = 16'hc088;
    LUT4 i14910_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14910_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_508 (.A(\select[4] ), .B(n29234), .C(n31503), .D(\read_size[2]_adj_314 ), 
         .Z(n9)) /* synthesis lut_function=(A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_508.init = 16'h8a88;
    LUT4 i14911_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14911_4_lut.init = 16'hc088;
    LUT4 i14912_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14912_4_lut.init = 16'hc088;
    LUT4 i14913_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14913_4_lut.init = 16'hc088;
    LUT4 i14914_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14914_4_lut.init = 16'hc088;
    LUT4 i2_4_lut_4_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(steps_reg[31]), .D(div_factor_reg[31]), .Z(n27420)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i2_4_lut_4_lut.init = 16'ha280;
    FD1S3IX steps_reg__i24 (.D(n4007[24]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4007[23]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4007[22]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4007[21]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4007[20]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4007[19]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4007[18]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4007[17]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4007[16]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4007[15]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4007[14]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4007[13]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4007[12]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4007[11]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4007[10]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4007[9]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4007[8]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4007[7]), .CK(debug_c_c), .CD(n31511), 
            .Q(\steps_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4007[6]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4007[5]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4007[4]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4007[3]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4007[2]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4007[1]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    PFUMX i22209 (.BLUT(n29767), .ALUT(n29768), .C0(\register_addr[0] ), 
          .Z(n29769));
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n31419), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n14522), .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n31419), .PD(n31511), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n14522), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n31419), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n31419), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n31419), .CD(n11208), 
            .CK(debug_c_c), .Q(control_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n14546), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n14546), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9304), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9304), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9304), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9304), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9304), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9304), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9304), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9304), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i13171_3_lut (.A(control_reg[7]), .B(div_factor_reg[7]), .C(\register_addr[1] ), 
         .Z(n19928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i13171_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_447 (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .Z(n31590)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut_rep_447.init = 16'heeee;
    LUT4 i2_2_lut_rep_397_3_lut_4_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(\register_addr[3] ), .D(\register_addr[2] ), .Z(n31540)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i2_2_lut_rep_397_3_lut_4_lut.init = 16'hfffe;
    LUT4 equal_66_i8_1_lut_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(\register_addr[3] ), .D(\register_addr[2] ), .Z(n6)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam equal_66_i8_1_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    PFUMX i22158 (.BLUT(n29716), .ALUT(n29717), .C0(\register_addr[1] ), 
          .Z(n29718));
    LUT4 mux_1575_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4006), 
         .Z(n4007[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4006), 
         .Z(n4007[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4006), 
         .Z(n4007[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4006), 
         .Z(n4007[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4006), 
         .Z(n4007[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4006), 
         .Z(n4007[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4006), 
         .Z(n4007[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4006), 
         .Z(n4007[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4006), 
         .Z(n4007[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4006), 
         .Z(n4007[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4006), 
         .Z(n4007[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4006), 
         .Z(n4007[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4006), 
         .Z(n4007[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4006), 
         .Z(n4007[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4006), 
         .Z(n4007[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4006), .Z(n4007[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4006), .Z(n4007[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4006), .Z(n4007[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4006), .Z(n4007[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4006), .Z(n4007[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4006), .Z(n4007[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4006), .Z(n4007[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4006), .Z(n4007[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4006), .Z(n4007[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i2_3_lut.init = 16'hcaca;
    LUT4 i14926_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8643[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14926_2_lut.init = 16'h2222;
    FD1P3AX read_value__i31 (.D(n27420), .SP(n2846), .CK(debug_c_c), .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1975_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7056[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1975_i4_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n31417), .SP(n10), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1575_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4006), .Z(n4007[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i1_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n14546), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=608, LSE_RLINE=621 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    LUT4 i14925_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8643[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14925_2_lut.init = 16'h2222;
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 mux_1975_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7056[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1975_i5_3_lut.init = 16'hcaca;
    LUT4 i14924_2_lut (.A(Stepper_Z_Dir_c), .B(\register_addr[0] ), .Z(n8643[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14924_2_lut.init = 16'h2222;
    LUT4 i22207_3_lut (.A(Stepper_Z_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n29767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22207_3_lut.init = 16'hcaca;
    LUT4 mux_1975_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7056[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1975_i6_3_lut.init = 16'hcaca;
    LUT4 i22208_3_lut (.A(n19910), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n29768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22208_3_lut.init = 16'hcaca;
    LUT4 i14923_2_lut (.A(Stepper_Z_En_c), .B(\register_addr[0] ), .Z(n8643[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14923_2_lut.init = 16'h2222;
    LUT4 mux_1975_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7056[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1975_i7_3_lut.init = 16'hcaca;
    PFUMX i13173 (.BLUT(n19928), .ALUT(n11), .C0(\register_addr[0] ), 
          .Z(n19930));
    LUT4 mux_1575_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4006), 
         .Z(n4007[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4006), 
         .Z(n4007[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4006), 
         .Z(n4007[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4006), 
         .Z(n4007[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4006), 
         .Z(n4007[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4006), 
         .Z(n4007[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1575_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4006), 
         .Z(n4007[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1575_i26_3_lut.init = 16'hcaca;
    PFUMX mux_1979_i4 (.BLUT(n8643[3]), .ALUT(n7056[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_1979_i5 (.BLUT(n8643[4]), .ALUT(n7056[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1979_i6 (.BLUT(n8643[5]), .ALUT(n7056[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1979_i7 (.BLUT(n8643[6]), .ALUT(n7056[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26850), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26849), .COUT(n26850), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26848), .COUT(n26849), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    PFUMX i22983 (.BLUT(n31614), .ALUT(n31615), .C0(\register_addr[0] ), 
          .Z(n31616));
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26847), .COUT(n26848), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26846), .COUT(n26847), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    ClockDivider step_clk_gen (.prev_step_clk(prev_step_clk), .n19910(n19910), 
            .step_clk(step_clk), .n31417(n31417), .n31511(n31511), .n10(n10), 
            .debug_c_c(debug_c_c), .n31410(n31410), .GND_net(GND_net), 
            .n16841(n16841), .div_factor_reg({div_factor_reg}), .n8263(n8263), 
            .n8297(n8297)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (prev_step_clk, n19910, step_clk, n31417, n31511, 
            n10, debug_c_c, n31410, GND_net, n16841, div_factor_reg, 
            n8263, n8297) /* synthesis syn_module_defined=1 */ ;
    input prev_step_clk;
    input n19910;
    output step_clk;
    output n31417;
    input n31511;
    output n10;
    input debug_c_c;
    input n31410;
    input GND_net;
    input n16841;
    input [31:0]div_factor_reg;
    output n8263;
    output n8297;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n8228;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n26602, n26601;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26600, n26599, n26598, n26597, n26596, n26595, n26594, 
        n26593, n26592, n26591, n26590, n26589, n26588, n26587, 
        n26786;
    wire [31:0]n40;
    
    wire n26785, n26586, n26585, n26584, n26583, n26922, n26921, 
        n26784, n26582, n26581, n26783, n26782, n26920, n26580, 
        n26919, n26918, n26917, n26781, n26916, n26915, n26914, 
        n26913, n26780, n26579, n26779, n26912, n26578, n26911, 
        n26577, n26910, n26576, n26778, n26777, n26909, n26776, 
        n26908, n26907, n26775, n26774, n26575, n26574, n26773, 
        n26573, n26772, n26572, n26571, n26771, n26570, n26569, 
        n26568, n26567, n26566, n26565, n26564, n26563, n26562, 
        n26561, n26560, n26559, n26558, n26557, n26556, n26555;
    
    LUT4 i2_3_lut_rep_274 (.A(prev_step_clk), .B(n19910), .C(step_clk), 
         .Z(n31417)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i2_3_lut_rep_274.init = 16'h4040;
    LUT4 i1_4_lut_4_lut (.A(prev_step_clk), .B(n19910), .C(step_clk), 
         .D(n31511), .Z(n10)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i1_4_lut_4_lut.init = 16'h004a;
    FD1S3IX clk_o_22 (.D(n8228), .CK(debug_c_c), .CD(n31511), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2675__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i0.GSR = "ENABLED";
    CCU2D sub_2073_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26602), .S1(n8228));
    defparam sub_2073_add_2_33.INIT0 = 16'h5555;
    defparam sub_2073_add_2_33.INIT1 = 16'h0000;
    defparam sub_2073_add_2_33.INJECT1_0 = "NO";
    defparam sub_2073_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26601), .COUT(n26602));
    defparam sub_2073_add_2_31.INIT0 = 16'h5999;
    defparam sub_2073_add_2_31.INIT1 = 16'h5999;
    defparam sub_2073_add_2_31.INJECT1_0 = "NO";
    defparam sub_2073_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26600), .COUT(n26601));
    defparam sub_2073_add_2_29.INIT0 = 16'h5999;
    defparam sub_2073_add_2_29.INIT1 = 16'h5999;
    defparam sub_2073_add_2_29.INJECT1_0 = "NO";
    defparam sub_2073_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26599), .COUT(n26600));
    defparam sub_2073_add_2_27.INIT0 = 16'h5999;
    defparam sub_2073_add_2_27.INIT1 = 16'h5999;
    defparam sub_2073_add_2_27.INJECT1_0 = "NO";
    defparam sub_2073_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26598), .COUT(n26599));
    defparam sub_2073_add_2_25.INIT0 = 16'h5999;
    defparam sub_2073_add_2_25.INIT1 = 16'h5999;
    defparam sub_2073_add_2_25.INJECT1_0 = "NO";
    defparam sub_2073_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26597), .COUT(n26598));
    defparam sub_2073_add_2_23.INIT0 = 16'h5999;
    defparam sub_2073_add_2_23.INIT1 = 16'h5999;
    defparam sub_2073_add_2_23.INJECT1_0 = "NO";
    defparam sub_2073_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26596), .COUT(n26597));
    defparam sub_2073_add_2_21.INIT0 = 16'h5999;
    defparam sub_2073_add_2_21.INIT1 = 16'h5999;
    defparam sub_2073_add_2_21.INJECT1_0 = "NO";
    defparam sub_2073_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26595), .COUT(n26596));
    defparam sub_2073_add_2_19.INIT0 = 16'h5999;
    defparam sub_2073_add_2_19.INIT1 = 16'h5999;
    defparam sub_2073_add_2_19.INJECT1_0 = "NO";
    defparam sub_2073_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26594), .COUT(n26595));
    defparam sub_2073_add_2_17.INIT0 = 16'h5999;
    defparam sub_2073_add_2_17.INIT1 = 16'h5999;
    defparam sub_2073_add_2_17.INJECT1_0 = "NO";
    defparam sub_2073_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26593), .COUT(n26594));
    defparam sub_2073_add_2_15.INIT0 = 16'h5999;
    defparam sub_2073_add_2_15.INIT1 = 16'h5999;
    defparam sub_2073_add_2_15.INJECT1_0 = "NO";
    defparam sub_2073_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26592), .COUT(n26593));
    defparam sub_2073_add_2_13.INIT0 = 16'h5999;
    defparam sub_2073_add_2_13.INIT1 = 16'h5999;
    defparam sub_2073_add_2_13.INJECT1_0 = "NO";
    defparam sub_2073_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26591), .COUT(n26592));
    defparam sub_2073_add_2_11.INIT0 = 16'h5999;
    defparam sub_2073_add_2_11.INIT1 = 16'h5999;
    defparam sub_2073_add_2_11.INJECT1_0 = "NO";
    defparam sub_2073_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26590), .COUT(n26591));
    defparam sub_2073_add_2_9.INIT0 = 16'h5999;
    defparam sub_2073_add_2_9.INIT1 = 16'h5999;
    defparam sub_2073_add_2_9.INJECT1_0 = "NO";
    defparam sub_2073_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26589), .COUT(n26590));
    defparam sub_2073_add_2_7.INIT0 = 16'h5999;
    defparam sub_2073_add_2_7.INIT1 = 16'h5999;
    defparam sub_2073_add_2_7.INJECT1_0 = "NO";
    defparam sub_2073_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2073_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26588), .COUT(n26589));
    defparam sub_2073_add_2_5.INIT0 = 16'h5999;
    defparam sub_2073_add_2_5.INIT1 = 16'h5999;
    defparam sub_2073_add_2_5.INJECT1_0 = "NO";
    defparam sub_2073_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26587), .COUT(n26588));
    defparam sub_2073_add_2_3.INIT0 = 16'h5999;
    defparam sub_2073_add_2_3.INIT1 = 16'h5999;
    defparam sub_2073_add_2_3.INJECT1_0 = "NO";
    defparam sub_2073_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26786), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26785), .COUT(n26786), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2073_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26587));
    defparam sub_2073_add_2_1.INIT0 = 16'h0000;
    defparam sub_2073_add_2_1.INIT1 = 16'h5999;
    defparam sub_2073_add_2_1.INJECT1_0 = "NO";
    defparam sub_2073_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26586), .S1(n8263));
    defparam sub_2075_add_2_33.INIT0 = 16'h5999;
    defparam sub_2075_add_2_33.INIT1 = 16'h0000;
    defparam sub_2075_add_2_33.INJECT1_0 = "NO";
    defparam sub_2075_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26585), .COUT(n26586));
    defparam sub_2075_add_2_31.INIT0 = 16'h5999;
    defparam sub_2075_add_2_31.INIT1 = 16'h5999;
    defparam sub_2075_add_2_31.INJECT1_0 = "NO";
    defparam sub_2075_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26584), .COUT(n26585));
    defparam sub_2075_add_2_29.INIT0 = 16'h5999;
    defparam sub_2075_add_2_29.INIT1 = 16'h5999;
    defparam sub_2075_add_2_29.INJECT1_0 = "NO";
    defparam sub_2075_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26583), .COUT(n26584));
    defparam sub_2075_add_2_27.INIT0 = 16'h5999;
    defparam sub_2075_add_2_27.INIT1 = 16'h5999;
    defparam sub_2075_add_2_27.INJECT1_0 = "NO";
    defparam sub_2075_add_2_27.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26922), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_33.INIT1 = 16'h0000;
    defparam count_2675_add_4_33.INJECT1_0 = "NO";
    defparam count_2675_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26921), .COUT(n26922), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_31.INJECT1_0 = "NO";
    defparam count_2675_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26784), .COUT(n26785), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26582), .COUT(n26583));
    defparam sub_2075_add_2_25.INIT0 = 16'h5999;
    defparam sub_2075_add_2_25.INIT1 = 16'h5999;
    defparam sub_2075_add_2_25.INJECT1_0 = "NO";
    defparam sub_2075_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26581), .COUT(n26582));
    defparam sub_2075_add_2_23.INIT0 = 16'h5999;
    defparam sub_2075_add_2_23.INIT1 = 16'h5999;
    defparam sub_2075_add_2_23.INJECT1_0 = "NO";
    defparam sub_2075_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26783), .COUT(n26784), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26782), .COUT(n26783), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26920), .COUT(n26921), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_29.INJECT1_0 = "NO";
    defparam count_2675_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26580), .COUT(n26581));
    defparam sub_2075_add_2_21.INIT0 = 16'h5999;
    defparam sub_2075_add_2_21.INIT1 = 16'h5999;
    defparam sub_2075_add_2_21.INJECT1_0 = "NO";
    defparam sub_2075_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26919), .COUT(n26920), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_27.INJECT1_0 = "NO";
    defparam count_2675_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26918), .COUT(n26919), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_25.INJECT1_0 = "NO";
    defparam count_2675_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26917), .COUT(n26918), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_23.INJECT1_0 = "NO";
    defparam count_2675_add_4_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26781), .COUT(n26782), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26916), .COUT(n26917), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_21.INJECT1_0 = "NO";
    defparam count_2675_add_4_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    CCU2D count_2675_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26915), .COUT(n26916), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_19.INJECT1_0 = "NO";
    defparam count_2675_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26914), .COUT(n26915), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_17.INJECT1_0 = "NO";
    defparam count_2675_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26913), .COUT(n26914), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_15.INJECT1_0 = "NO";
    defparam count_2675_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26780), .COUT(n26781), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    CCU2D sub_2075_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26579), .COUT(n26580));
    defparam sub_2075_add_2_19.INIT0 = 16'h5999;
    defparam sub_2075_add_2_19.INIT1 = 16'h5999;
    defparam sub_2075_add_2_19.INJECT1_0 = "NO";
    defparam sub_2075_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26779), .COUT(n26780), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26912), .COUT(n26913), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_13.INJECT1_0 = "NO";
    defparam count_2675_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26578), .COUT(n26579));
    defparam sub_2075_add_2_17.INIT0 = 16'h5999;
    defparam sub_2075_add_2_17.INIT1 = 16'h5999;
    defparam sub_2075_add_2_17.INJECT1_0 = "NO";
    defparam sub_2075_add_2_17.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    CCU2D count_2675_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26911), .COUT(n26912), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_11.INJECT1_0 = "NO";
    defparam count_2675_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26577), .COUT(n26578));
    defparam sub_2075_add_2_15.INIT0 = 16'h5999;
    defparam sub_2075_add_2_15.INIT1 = 16'h5999;
    defparam sub_2075_add_2_15.INJECT1_0 = "NO";
    defparam sub_2075_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26910), .COUT(n26911), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_9.INJECT1_0 = "NO";
    defparam count_2675_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26576), .COUT(n26577));
    defparam sub_2075_add_2_13.INIT0 = 16'h5999;
    defparam sub_2075_add_2_13.INIT1 = 16'h5999;
    defparam sub_2075_add_2_13.INJECT1_0 = "NO";
    defparam sub_2075_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26778), .COUT(n26779), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26777), .COUT(n26778), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26909), .COUT(n26910), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_7.INJECT1_0 = "NO";
    defparam count_2675_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26776), .COUT(n26777), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26908), .COUT(n26909), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_5.INJECT1_0 = "NO";
    defparam count_2675_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26907), .COUT(n26908), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_3.INJECT1_0 = "NO";
    defparam count_2675_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26775), .COUT(n26776), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26907), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_1.INIT0 = 16'hF000;
    defparam count_2675_add_4_1.INIT1 = 16'h0555;
    defparam count_2675_add_4_1.INJECT1_0 = "NO";
    defparam count_2675_add_4_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26774), .COUT(n26775), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26575), .COUT(n26576));
    defparam sub_2075_add_2_11.INIT0 = 16'h5999;
    defparam sub_2075_add_2_11.INIT1 = 16'h5999;
    defparam sub_2075_add_2_11.INJECT1_0 = "NO";
    defparam sub_2075_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26574), .COUT(n26575));
    defparam sub_2075_add_2_9.INIT0 = 16'h5999;
    defparam sub_2075_add_2_9.INIT1 = 16'h5999;
    defparam sub_2075_add_2_9.INJECT1_0 = "NO";
    defparam sub_2075_add_2_9.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26773), .COUT(n26774), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31410), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31410), .PD(n16841), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2075_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26573), .COUT(n26574));
    defparam sub_2075_add_2_7.INIT0 = 16'h5999;
    defparam sub_2075_add_2_7.INIT1 = 16'h5999;
    defparam sub_2075_add_2_7.INJECT1_0 = "NO";
    defparam sub_2075_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26772), .COUT(n26773), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    FD1S3IX count_2675__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i1.GSR = "ENABLED";
    CCU2D sub_2075_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26572), .COUT(n26573));
    defparam sub_2075_add_2_5.INIT0 = 16'h5999;
    defparam sub_2075_add_2_5.INIT1 = 16'h5999;
    defparam sub_2075_add_2_5.INJECT1_0 = "NO";
    defparam sub_2075_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26571), .COUT(n26572));
    defparam sub_2075_add_2_3.INIT0 = 16'h5999;
    defparam sub_2075_add_2_3.INIT1 = 16'h5999;
    defparam sub_2075_add_2_3.INJECT1_0 = "NO";
    defparam sub_2075_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2075_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26571));
    defparam sub_2075_add_2_1.INIT0 = 16'h0000;
    defparam sub_2075_add_2_1.INIT1 = 16'h5999;
    defparam sub_2075_add_2_1.INJECT1_0 = "NO";
    defparam sub_2075_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26771), .COUT(n26772), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26570), .S1(n8297));
    defparam sub_2076_add_2_33.INIT0 = 16'hf555;
    defparam sub_2076_add_2_33.INIT1 = 16'h0000;
    defparam sub_2076_add_2_33.INJECT1_0 = "NO";
    defparam sub_2076_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26771), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26569), .COUT(n26570));
    defparam sub_2076_add_2_31.INIT0 = 16'hf555;
    defparam sub_2076_add_2_31.INIT1 = 16'hf555;
    defparam sub_2076_add_2_31.INJECT1_0 = "NO";
    defparam sub_2076_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26568), .COUT(n26569));
    defparam sub_2076_add_2_29.INIT0 = 16'hf555;
    defparam sub_2076_add_2_29.INIT1 = 16'hf555;
    defparam sub_2076_add_2_29.INJECT1_0 = "NO";
    defparam sub_2076_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26567), .COUT(n26568));
    defparam sub_2076_add_2_27.INIT0 = 16'hf555;
    defparam sub_2076_add_2_27.INIT1 = 16'hf555;
    defparam sub_2076_add_2_27.INJECT1_0 = "NO";
    defparam sub_2076_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26566), .COUT(n26567));
    defparam sub_2076_add_2_25.INIT0 = 16'hf555;
    defparam sub_2076_add_2_25.INIT1 = 16'hf555;
    defparam sub_2076_add_2_25.INJECT1_0 = "NO";
    defparam sub_2076_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26565), .COUT(n26566));
    defparam sub_2076_add_2_23.INIT0 = 16'hf555;
    defparam sub_2076_add_2_23.INIT1 = 16'hf555;
    defparam sub_2076_add_2_23.INJECT1_0 = "NO";
    defparam sub_2076_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26564), .COUT(n26565));
    defparam sub_2076_add_2_21.INIT0 = 16'hf555;
    defparam sub_2076_add_2_21.INIT1 = 16'hf555;
    defparam sub_2076_add_2_21.INJECT1_0 = "NO";
    defparam sub_2076_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26563), .COUT(n26564));
    defparam sub_2076_add_2_19.INIT0 = 16'hf555;
    defparam sub_2076_add_2_19.INIT1 = 16'hf555;
    defparam sub_2076_add_2_19.INJECT1_0 = "NO";
    defparam sub_2076_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26562), .COUT(n26563));
    defparam sub_2076_add_2_17.INIT0 = 16'hf555;
    defparam sub_2076_add_2_17.INIT1 = 16'hf555;
    defparam sub_2076_add_2_17.INJECT1_0 = "NO";
    defparam sub_2076_add_2_17.INJECT1_1 = "NO";
    FD1S3IX count_2675__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i2.GSR = "ENABLED";
    FD1S3IX count_2675__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i3.GSR = "ENABLED";
    FD1S3IX count_2675__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i4.GSR = "ENABLED";
    FD1S3IX count_2675__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i5.GSR = "ENABLED";
    FD1S3IX count_2675__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i6.GSR = "ENABLED";
    FD1S3IX count_2675__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i7.GSR = "ENABLED";
    FD1S3IX count_2675__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i8.GSR = "ENABLED";
    FD1S3IX count_2675__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i9.GSR = "ENABLED";
    FD1S3IX count_2675__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i10.GSR = "ENABLED";
    FD1S3IX count_2675__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i11.GSR = "ENABLED";
    FD1S3IX count_2675__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i12.GSR = "ENABLED";
    FD1S3IX count_2675__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i13.GSR = "ENABLED";
    FD1S3IX count_2675__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i14.GSR = "ENABLED";
    FD1S3IX count_2675__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i15.GSR = "ENABLED";
    FD1S3IX count_2675__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i16.GSR = "ENABLED";
    FD1S3IX count_2675__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i17.GSR = "ENABLED";
    FD1S3IX count_2675__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i18.GSR = "ENABLED";
    FD1S3IX count_2675__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i19.GSR = "ENABLED";
    FD1S3IX count_2675__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i20.GSR = "ENABLED";
    FD1S3IX count_2675__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i21.GSR = "ENABLED";
    FD1S3IX count_2675__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i22.GSR = "ENABLED";
    FD1S3IX count_2675__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i23.GSR = "ENABLED";
    FD1S3IX count_2675__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i24.GSR = "ENABLED";
    FD1S3IX count_2675__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i25.GSR = "ENABLED";
    FD1S3IX count_2675__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i26.GSR = "ENABLED";
    FD1S3IX count_2675__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i27.GSR = "ENABLED";
    FD1S3IX count_2675__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i28.GSR = "ENABLED";
    FD1S3IX count_2675__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i29.GSR = "ENABLED";
    FD1S3IX count_2675__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i30.GSR = "ENABLED";
    FD1S3IX count_2675__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i31.GSR = "ENABLED";
    CCU2D sub_2076_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26561), .COUT(n26562));
    defparam sub_2076_add_2_15.INIT0 = 16'hf555;
    defparam sub_2076_add_2_15.INIT1 = 16'hf555;
    defparam sub_2076_add_2_15.INJECT1_0 = "NO";
    defparam sub_2076_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26560), .COUT(n26561));
    defparam sub_2076_add_2_13.INIT0 = 16'hf555;
    defparam sub_2076_add_2_13.INIT1 = 16'hf555;
    defparam sub_2076_add_2_13.INJECT1_0 = "NO";
    defparam sub_2076_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26559), .COUT(n26560));
    defparam sub_2076_add_2_11.INIT0 = 16'hf555;
    defparam sub_2076_add_2_11.INIT1 = 16'hf555;
    defparam sub_2076_add_2_11.INJECT1_0 = "NO";
    defparam sub_2076_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26558), .COUT(n26559));
    defparam sub_2076_add_2_9.INIT0 = 16'hf555;
    defparam sub_2076_add_2_9.INIT1 = 16'hf555;
    defparam sub_2076_add_2_9.INJECT1_0 = "NO";
    defparam sub_2076_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26557), .COUT(n26558));
    defparam sub_2076_add_2_7.INIT0 = 16'hf555;
    defparam sub_2076_add_2_7.INIT1 = 16'hf555;
    defparam sub_2076_add_2_7.INJECT1_0 = "NO";
    defparam sub_2076_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26556), .COUT(n26557));
    defparam sub_2076_add_2_5.INIT0 = 16'hf555;
    defparam sub_2076_add_2_5.INIT1 = 16'hf555;
    defparam sub_2076_add_2_5.INJECT1_0 = "NO";
    defparam sub_2076_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26555), .COUT(n26556));
    defparam sub_2076_add_2_3.INIT0 = 16'hf555;
    defparam sub_2076_add_2_3.INIT1 = 16'hf555;
    defparam sub_2076_add_2_3.INJECT1_0 = "NO";
    defparam sub_2076_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26555));
    defparam sub_2076_add_2_1.INIT0 = 16'h0000;
    defparam sub_2076_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2076_add_2_1.INJECT1_0 = "NO";
    defparam sub_2076_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (debug_c_c, VCC_net, GND_net, 
            Stepper_Y_nFault_c, n31511, n4094, \read_size[0] , n14650, 
            n27751, Stepper_Y_M0_c_0, databus, prev_step_clk, step_clk, 
            limit_latched, prev_limit_latched, n9300, prev_select, n31445, 
            n29270, n29491, Stepper_Y_M1_c_1, \register_addr[0] , \div_factor_reg[9] , 
            \div_factor_reg[6] , \div_factor_reg[5] , \div_factor_reg[4] , 
            \div_factor_reg[3] , \control_reg[7] , n12148, Stepper_Y_En_c, 
            Stepper_Y_Dir_c, \control_reg[4] , \control_reg[3] , Stepper_Y_M2_c_2, 
            \read_size[2] , n29199, \steps_reg[9] , \steps_reg[6] , 
            \steps_reg[5] , \steps_reg[4] , \steps_reg[3] , read_value, 
            n9547, \register_addr[1] , n29112, limit_c_1, int_step, 
            n22, n31418, n29113, n21213, n21221, n28826, n6807, 
            n32, n27483, n224, n8635, n8193, n31407, n16840, n8159) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    input n31511;
    input [31:0]n4094;
    output \read_size[0] ;
    input n14650;
    input n27751;
    output Stepper_Y_M0_c_0;
    input [31:0]databus;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    input n9300;
    output prev_select;
    input n31445;
    input n29270;
    input n29491;
    output Stepper_Y_M1_c_1;
    input \register_addr[0] ;
    output \div_factor_reg[9] ;
    output \div_factor_reg[6] ;
    output \div_factor_reg[5] ;
    output \div_factor_reg[4] ;
    output \div_factor_reg[3] ;
    output \control_reg[7] ;
    input n12148;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output \control_reg[4] ;
    output \control_reg[3] ;
    output Stepper_Y_M2_c_2;
    output \read_size[2] ;
    input n29199;
    output \steps_reg[9] ;
    output \steps_reg[6] ;
    output \steps_reg[5] ;
    output \steps_reg[4] ;
    output \steps_reg[3] ;
    output [31:0]read_value;
    input n9547;
    input \register_addr[1] ;
    input n29112;
    input limit_c_1;
    output int_step;
    input n22;
    input n31418;
    input n29113;
    input n21213;
    input n21221;
    input n28826;
    input n6807;
    input n32;
    output n27483;
    output [31:0]n224;
    input n8635;
    output n8193;
    input n31407;
    input n16840;
    output n8159;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire fault_latched;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n13923, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n29713, n29714, n29740, n29741, n29742;
    wire [31:0]n100;
    
    wire n29686, n29687, n29688, n29715;
    wire [31:0]n6742;
    
    wire n29132, n29120, n29133, n29134, n29135, n29131, n29130, 
        n29129, n29128, n29125, n29127, n29126, n29124, n29123, 
        n29122, n29121, n29114, n29118, n29116, n29119, n29117, 
        n29115;
    wire [31:0]n6778;
    
    wire n49, n62, n58, n50, n41, n60, n54, n42, n52, n38, 
        n56, n46, n26866, n26865, n26864, n26863, n26862, n26861, 
        n26860, n26859, n26858, n26857, n26856, n26855, n26854, 
        n26853, n26852, n26851;
    
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4094[0]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n27751), .SP(n14650), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n13923), .CD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31445), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31445), .B(prev_select), .C(n29270), 
         .D(n29491), .Z(n13923)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i22153_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22153_3_lut.init = 16'hcaca;
    LUT4 i22154_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22154_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9300), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9300), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9300), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9300), .PD(n31511), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9300), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9300), .PD(n31511), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9300), .PD(n31511), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(\div_factor_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n9300), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13923), .CD(n12148), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13923), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13923), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13923), .CD(n31511), 
            .CK(debug_c_c), .Q(\control_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13923), .PD(n31511), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13923), .CD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13923), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    PFUMX i22182 (.BLUT(n29740), .ALUT(n29741), .C0(\register_addr[0] ), 
          .Z(n29742));
    FD1P3AX read_size__i2 (.D(n29199), .SP(n14650), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n4094[31]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4094[30]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4094[29]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4094[28]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4094[27]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4094[26]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4094[25]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4094[24]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4094[23]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4094[22]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4094[21]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4094[20]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4094[19]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4094[18]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4094[17]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4094[16]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4094[15]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4094[14]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4094[13]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4094[12]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4094[11]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4094[10]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4094[9]), .CK(debug_c_c), .CD(n31511), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4094[8]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4094[7]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4094[6]), .CK(debug_c_c), .CD(n31511), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4094[5]), .CK(debug_c_c), .CD(n31511), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4094[4]), .CK(debug_c_c), .CD(n31511), 
            .Q(\steps_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4094[3]), .CK(debug_c_c), .CD(n31511), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4094[2]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4094[1]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    PFUMX i22128 (.BLUT(n29686), .ALUT(n29687), .C0(\register_addr[1] ), 
          .Z(n29688));
    PFUMX i22155 (.BLUT(n29713), .ALUT(n29714), .C0(\register_addr[1] ), 
          .Z(n29715));
    LUT4 i22126_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n29686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22126_3_lut.init = 16'hcaca;
    LUT4 i22127_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n29687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22127_3_lut.init = 16'hcaca;
    LUT4 mux_1949_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6742[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1949_i8_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i30 (.D(n29132), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29120), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29133), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29134), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29135), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29131), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29130), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29129), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29128), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29125), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29127), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29126), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29124), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29123), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29122), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29121), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(div_factor_reg[30]), .B(n29112), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29132)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_483 (.A(div_factor_reg[29]), .B(n29112), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29120)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_483.init = 16'hc088;
    FD1P3AX int_step_182 (.D(n31418), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29114), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29118), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29116), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29119), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29117), .SP(n14650), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29113), .SP(n14650), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29115), .SP(n14650), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6778[7]), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n21213), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n21221), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n28826), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6807), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29742), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29715), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_484 (.A(div_factor_reg[28]), .B(n29112), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n29133)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_484.init = 16'hc088;
    LUT4 i1_4_lut_adj_485 (.A(div_factor_reg[27]), .B(n29112), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n29134)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_485.init = 16'hc088;
    LUT4 i1_4_lut_adj_486 (.A(div_factor_reg[26]), .B(n29112), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n29135)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_486.init = 16'hc088;
    LUT4 i1_4_lut_adj_487 (.A(div_factor_reg[25]), .B(n29112), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n29131)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_487.init = 16'hc088;
    LUT4 i1_4_lut_adj_488 (.A(div_factor_reg[24]), .B(n29112), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n29130)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_488.init = 16'hc088;
    LUT4 i1_4_lut_adj_489 (.A(div_factor_reg[23]), .B(n29112), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n29129)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_489.init = 16'hc088;
    LUT4 i1_4_lut_adj_490 (.A(div_factor_reg[22]), .B(n29112), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n29128)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_490.init = 16'hc088;
    LUT4 i22180_3_lut (.A(Stepper_Y_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n29740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22180_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n29688), .SP(n14650), .CD(n9547), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=593, LSE_RLINE=606 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i22181_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n29741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22181_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_491 (.A(div_factor_reg[21]), .B(n29112), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n29125)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_491.init = 16'hc088;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27483)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_492 (.A(div_factor_reg[20]), .B(n29112), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n29127)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_492.init = 16'hc088;
    LUT4 i1_4_lut_adj_493 (.A(div_factor_reg[19]), .B(n29112), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n29126)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_493.init = 16'hc088;
    LUT4 i1_4_lut_adj_494 (.A(div_factor_reg[18]), .B(n29112), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n29124)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_494.init = 16'hc088;
    LUT4 i1_4_lut_adj_495 (.A(div_factor_reg[17]), .B(n29112), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n29123)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_495.init = 16'hc088;
    LUT4 i1_4_lut_adj_496 (.A(div_factor_reg[16]), .B(n29112), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n29122)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_496.init = 16'hc088;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_497 (.A(div_factor_reg[15]), .B(n29112), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n29121)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_497.init = 16'hc088;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(\steps_reg[4] ), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_498 (.A(div_factor_reg[14]), .B(n29112), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n29114)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_498.init = 16'hc088;
    LUT4 i1_4_lut_adj_499 (.A(div_factor_reg[13]), .B(n29112), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n29118)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_499.init = 16'hc088;
    LUT4 i1_4_lut_adj_500 (.A(div_factor_reg[12]), .B(n29112), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n29116)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_500.init = 16'hc088;
    LUT4 i1_4_lut_adj_501 (.A(div_factor_reg[11]), .B(n29112), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n29119)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_501.init = 16'hc088;
    LUT4 i1_4_lut_adj_502 (.A(div_factor_reg[10]), .B(n29112), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n29117)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_502.init = 16'hc088;
    LUT4 i1_4_lut_adj_503 (.A(div_factor_reg[8]), .B(n29112), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29115)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_503.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26866), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26865), .COUT(n26866), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26864), .COUT(n26865), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26863), .COUT(n26864), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26862), .COUT(n26863), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26861), .COUT(n26862), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26860), .COUT(n26861), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26859), .COUT(n26860), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26858), .COUT(n26859), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26857), .COUT(n26858), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26856), .COUT(n26857), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26855), .COUT(n26856), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    PFUMX mux_1953_i8 (.BLUT(n8635), .ALUT(n6742[7]), .C0(\register_addr[1] ), 
          .Z(n6778[7]));
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26854), .COUT(n26855), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 i14927_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14927_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26853), .COUT(n26854), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26852), .COUT(n26853), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26851), .COUT(n26852), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n26851), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    ClockDivider_U7 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n31511(n31511), .div_factor_reg({div_factor_reg[31:10], 
            \div_factor_reg[9] , div_factor_reg[8:7], \div_factor_reg[6] , 
            \div_factor_reg[5] , \div_factor_reg[4] , \div_factor_reg[3] , 
            div_factor_reg[2:0]}), .n8193(n8193), .n31407(n31407), .n16840(n16840), 
            .n8159(n8159)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (GND_net, step_clk, debug_c_c, n31511, div_factor_reg, 
            n8193, n31407, n16840, n8159) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31511;
    input [31:0]div_factor_reg;
    output n8193;
    input n31407;
    input n16840;
    output n8159;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26628;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n40;
    
    wire n26629, n26627, n26626, n26625, n26624, n26623, n26622, 
        n26621, n8124, n26620, n26619, n26618, n26617, n26616, 
        n26615, n26614, n26613, n26612, n26611, n26610, n26609, 
        n26802;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26608, n26801;
    wire [31:0]n134;
    
    wire n26800, n26799, n26798, n26797, n26796, n26607, n26795, 
        n26794, n26606, n26605, n26793, n26604, n26603, n26792, 
        n26791, n26790, n26789, n26788, n26787, n26650, n26649, 
        n26648, n26647, n26646, n26645, n26644, n26643, n27034, 
        n26642, n27033, n27032, n27031, n27030, n27029, n27028, 
        n27027, n27026, n26641, n26640, n27025, n27024, n27023, 
        n26639, n27022, n26638, n27021, n27020, n27019, n26637, 
        n26636, n26635, n26634, n26633, n26632, n26631, n26630;
    
    CCU2D sub_2070_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26628), .COUT(n26629));
    defparam sub_2070_add_2_21.INIT0 = 16'h5999;
    defparam sub_2070_add_2_21.INIT1 = 16'h5999;
    defparam sub_2070_add_2_21.INJECT1_0 = "NO";
    defparam sub_2070_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26627), .COUT(n26628));
    defparam sub_2070_add_2_19.INIT0 = 16'h5999;
    defparam sub_2070_add_2_19.INIT1 = 16'h5999;
    defparam sub_2070_add_2_19.INJECT1_0 = "NO";
    defparam sub_2070_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26626), .COUT(n26627));
    defparam sub_2070_add_2_17.INIT0 = 16'h5999;
    defparam sub_2070_add_2_17.INIT1 = 16'h5999;
    defparam sub_2070_add_2_17.INJECT1_0 = "NO";
    defparam sub_2070_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26625), .COUT(n26626));
    defparam sub_2070_add_2_15.INIT0 = 16'h5999;
    defparam sub_2070_add_2_15.INIT1 = 16'h5999;
    defparam sub_2070_add_2_15.INJECT1_0 = "NO";
    defparam sub_2070_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26624), .COUT(n26625));
    defparam sub_2070_add_2_13.INIT0 = 16'h5999;
    defparam sub_2070_add_2_13.INIT1 = 16'h5999;
    defparam sub_2070_add_2_13.INJECT1_0 = "NO";
    defparam sub_2070_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26623), .COUT(n26624));
    defparam sub_2070_add_2_11.INIT0 = 16'h5999;
    defparam sub_2070_add_2_11.INIT1 = 16'h5999;
    defparam sub_2070_add_2_11.INJECT1_0 = "NO";
    defparam sub_2070_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26622), .COUT(n26623));
    defparam sub_2070_add_2_9.INIT0 = 16'h5999;
    defparam sub_2070_add_2_9.INIT1 = 16'h5999;
    defparam sub_2070_add_2_9.INJECT1_0 = "NO";
    defparam sub_2070_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26621), .COUT(n26622));
    defparam sub_2070_add_2_7.INIT0 = 16'h5999;
    defparam sub_2070_add_2_7.INIT1 = 16'h5999;
    defparam sub_2070_add_2_7.INJECT1_0 = "NO";
    defparam sub_2070_add_2_7.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8124), .CK(debug_c_c), .CD(n31511), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2070_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26620), .COUT(n26621));
    defparam sub_2070_add_2_5.INIT0 = 16'h5999;
    defparam sub_2070_add_2_5.INIT1 = 16'h5999;
    defparam sub_2070_add_2_5.INJECT1_0 = "NO";
    defparam sub_2070_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26619), .COUT(n26620));
    defparam sub_2070_add_2_3.INIT0 = 16'h5999;
    defparam sub_2070_add_2_3.INIT1 = 16'h5999;
    defparam sub_2070_add_2_3.INJECT1_0 = "NO";
    defparam sub_2070_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26619));
    defparam sub_2070_add_2_1.INIT0 = 16'h0000;
    defparam sub_2070_add_2_1.INIT1 = 16'h5999;
    defparam sub_2070_add_2_1.INJECT1_0 = "NO";
    defparam sub_2070_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26618), .S1(n8193));
    defparam sub_2071_add_2_33.INIT0 = 16'hf555;
    defparam sub_2071_add_2_33.INIT1 = 16'h0000;
    defparam sub_2071_add_2_33.INJECT1_0 = "NO";
    defparam sub_2071_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26617), .COUT(n26618));
    defparam sub_2071_add_2_31.INIT0 = 16'hf555;
    defparam sub_2071_add_2_31.INIT1 = 16'hf555;
    defparam sub_2071_add_2_31.INJECT1_0 = "NO";
    defparam sub_2071_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26616), .COUT(n26617));
    defparam sub_2071_add_2_29.INIT0 = 16'hf555;
    defparam sub_2071_add_2_29.INIT1 = 16'hf555;
    defparam sub_2071_add_2_29.INJECT1_0 = "NO";
    defparam sub_2071_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26615), .COUT(n26616));
    defparam sub_2071_add_2_27.INIT0 = 16'hf555;
    defparam sub_2071_add_2_27.INIT1 = 16'hf555;
    defparam sub_2071_add_2_27.INJECT1_0 = "NO";
    defparam sub_2071_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26614), .COUT(n26615));
    defparam sub_2071_add_2_25.INIT0 = 16'hf555;
    defparam sub_2071_add_2_25.INIT1 = 16'hf555;
    defparam sub_2071_add_2_25.INJECT1_0 = "NO";
    defparam sub_2071_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26613), .COUT(n26614));
    defparam sub_2071_add_2_23.INIT0 = 16'hf555;
    defparam sub_2071_add_2_23.INIT1 = 16'hf555;
    defparam sub_2071_add_2_23.INJECT1_0 = "NO";
    defparam sub_2071_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26612), .COUT(n26613));
    defparam sub_2071_add_2_21.INIT0 = 16'hf555;
    defparam sub_2071_add_2_21.INIT1 = 16'hf555;
    defparam sub_2071_add_2_21.INJECT1_0 = "NO";
    defparam sub_2071_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26611), .COUT(n26612));
    defparam sub_2071_add_2_19.INIT0 = 16'hf555;
    defparam sub_2071_add_2_19.INIT1 = 16'hf555;
    defparam sub_2071_add_2_19.INJECT1_0 = "NO";
    defparam sub_2071_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26610), .COUT(n26611));
    defparam sub_2071_add_2_17.INIT0 = 16'hf555;
    defparam sub_2071_add_2_17.INIT1 = 16'hf555;
    defparam sub_2071_add_2_17.INJECT1_0 = "NO";
    defparam sub_2071_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26609), .COUT(n26610));
    defparam sub_2071_add_2_15.INIT0 = 16'hf555;
    defparam sub_2071_add_2_15.INIT1 = 16'hf555;
    defparam sub_2071_add_2_15.INJECT1_0 = "NO";
    defparam sub_2071_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26802), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26608), .COUT(n26609));
    defparam sub_2071_add_2_13.INIT0 = 16'hf555;
    defparam sub_2071_add_2_13.INIT1 = 16'hf555;
    defparam sub_2071_add_2_13.INJECT1_0 = "NO";
    defparam sub_2071_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26801), .COUT(n26802), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    FD1S3IX count_2674__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26800), .COUT(n26801), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26799), .COUT(n26800), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26798), .COUT(n26799), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26797), .COUT(n26798), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26796), .COUT(n26797), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26607), .COUT(n26608));
    defparam sub_2071_add_2_11.INIT0 = 16'hf555;
    defparam sub_2071_add_2_11.INIT1 = 16'hf555;
    defparam sub_2071_add_2_11.INJECT1_0 = "NO";
    defparam sub_2071_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26795), .COUT(n26796), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26794), .COUT(n26795), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26606), .COUT(n26607));
    defparam sub_2071_add_2_9.INIT0 = 16'hf555;
    defparam sub_2071_add_2_9.INIT1 = 16'hf555;
    defparam sub_2071_add_2_9.INJECT1_0 = "NO";
    defparam sub_2071_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26605), .COUT(n26606));
    defparam sub_2071_add_2_7.INIT0 = 16'hf555;
    defparam sub_2071_add_2_7.INIT1 = 16'hf555;
    defparam sub_2071_add_2_7.INJECT1_0 = "NO";
    defparam sub_2071_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26793), .COUT(n26794), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26604), .COUT(n26605));
    defparam sub_2071_add_2_5.INIT0 = 16'hf555;
    defparam sub_2071_add_2_5.INIT1 = 16'hf555;
    defparam sub_2071_add_2_5.INJECT1_0 = "NO";
    defparam sub_2071_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26603), .COUT(n26604));
    defparam sub_2071_add_2_3.INIT0 = 16'hf555;
    defparam sub_2071_add_2_3.INIT1 = 16'hf555;
    defparam sub_2071_add_2_3.INJECT1_0 = "NO";
    defparam sub_2071_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26792), .COUT(n26793), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26603));
    defparam sub_2071_add_2_1.INIT0 = 16'h0000;
    defparam sub_2071_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2071_add_2_1.INJECT1_0 = "NO";
    defparam sub_2071_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26791), .COUT(n26792), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26790), .COUT(n26791), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26789), .COUT(n26790), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26788), .COUT(n26789), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26787), .COUT(n26788), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26787), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31407), .CD(n16840), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31407), .PD(n16840), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2068_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26650), .S1(n8124));
    defparam sub_2068_add_2_33.INIT0 = 16'h5555;
    defparam sub_2068_add_2_33.INIT1 = 16'h0000;
    defparam sub_2068_add_2_33.INJECT1_0 = "NO";
    defparam sub_2068_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26649), .COUT(n26650));
    defparam sub_2068_add_2_31.INIT0 = 16'h5999;
    defparam sub_2068_add_2_31.INIT1 = 16'h5999;
    defparam sub_2068_add_2_31.INJECT1_0 = "NO";
    defparam sub_2068_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26648), .COUT(n26649));
    defparam sub_2068_add_2_29.INIT0 = 16'h5999;
    defparam sub_2068_add_2_29.INIT1 = 16'h5999;
    defparam sub_2068_add_2_29.INJECT1_0 = "NO";
    defparam sub_2068_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26647), .COUT(n26648));
    defparam sub_2068_add_2_27.INIT0 = 16'h5999;
    defparam sub_2068_add_2_27.INIT1 = 16'h5999;
    defparam sub_2068_add_2_27.INJECT1_0 = "NO";
    defparam sub_2068_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26646), .COUT(n26647));
    defparam sub_2068_add_2_25.INIT0 = 16'h5999;
    defparam sub_2068_add_2_25.INIT1 = 16'h5999;
    defparam sub_2068_add_2_25.INJECT1_0 = "NO";
    defparam sub_2068_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26645), .COUT(n26646));
    defparam sub_2068_add_2_23.INIT0 = 16'h5999;
    defparam sub_2068_add_2_23.INIT1 = 16'h5999;
    defparam sub_2068_add_2_23.INJECT1_0 = "NO";
    defparam sub_2068_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26644), .COUT(n26645));
    defparam sub_2068_add_2_21.INIT0 = 16'h5999;
    defparam sub_2068_add_2_21.INIT1 = 16'h5999;
    defparam sub_2068_add_2_21.INJECT1_0 = "NO";
    defparam sub_2068_add_2_21.INJECT1_1 = "NO";
    FD1S3IX count_2674__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i1.GSR = "ENABLED";
    FD1S3IX count_2674__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i2.GSR = "ENABLED";
    FD1S3IX count_2674__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i3.GSR = "ENABLED";
    FD1S3IX count_2674__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i4.GSR = "ENABLED";
    FD1S3IX count_2674__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i5.GSR = "ENABLED";
    FD1S3IX count_2674__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i6.GSR = "ENABLED";
    FD1S3IX count_2674__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i7.GSR = "ENABLED";
    FD1S3IX count_2674__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i8.GSR = "ENABLED";
    FD1S3IX count_2674__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i9.GSR = "ENABLED";
    FD1S3IX count_2674__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i10.GSR = "ENABLED";
    FD1S3IX count_2674__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i11.GSR = "ENABLED";
    FD1S3IX count_2674__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i12.GSR = "ENABLED";
    FD1S3IX count_2674__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i13.GSR = "ENABLED";
    FD1S3IX count_2674__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i14.GSR = "ENABLED";
    FD1S3IX count_2674__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i15.GSR = "ENABLED";
    FD1S3IX count_2674__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i16.GSR = "ENABLED";
    FD1S3IX count_2674__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i17.GSR = "ENABLED";
    FD1S3IX count_2674__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i18.GSR = "ENABLED";
    FD1S3IX count_2674__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i19.GSR = "ENABLED";
    FD1S3IX count_2674__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i20.GSR = "ENABLED";
    FD1S3IX count_2674__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i21.GSR = "ENABLED";
    FD1S3IX count_2674__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i22.GSR = "ENABLED";
    FD1S3IX count_2674__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i23.GSR = "ENABLED";
    FD1S3IX count_2674__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i24.GSR = "ENABLED";
    FD1S3IX count_2674__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i25.GSR = "ENABLED";
    FD1S3IX count_2674__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i26.GSR = "ENABLED";
    FD1S3IX count_2674__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i27.GSR = "ENABLED";
    FD1S3IX count_2674__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i28.GSR = "ENABLED";
    FD1S3IX count_2674__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i29.GSR = "ENABLED";
    FD1S3IX count_2674__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i30.GSR = "ENABLED";
    FD1S3IX count_2674__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31407), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i31.GSR = "ENABLED";
    CCU2D sub_2068_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26643), .COUT(n26644));
    defparam sub_2068_add_2_19.INIT0 = 16'h5999;
    defparam sub_2068_add_2_19.INIT1 = 16'h5999;
    defparam sub_2068_add_2_19.INJECT1_0 = "NO";
    defparam sub_2068_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27034), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_33.INIT1 = 16'h0000;
    defparam count_2674_add_4_33.INJECT1_0 = "NO";
    defparam count_2674_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26642), .COUT(n26643));
    defparam sub_2068_add_2_17.INIT0 = 16'h5999;
    defparam sub_2068_add_2_17.INIT1 = 16'h5999;
    defparam sub_2068_add_2_17.INJECT1_0 = "NO";
    defparam sub_2068_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27033), .COUT(n27034), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_31.INJECT1_0 = "NO";
    defparam count_2674_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27032), .COUT(n27033), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_29.INJECT1_0 = "NO";
    defparam count_2674_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27031), .COUT(n27032), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_27.INJECT1_0 = "NO";
    defparam count_2674_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27030), .COUT(n27031), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_25.INJECT1_0 = "NO";
    defparam count_2674_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27029), .COUT(n27030), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_23.INJECT1_0 = "NO";
    defparam count_2674_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27028), .COUT(n27029), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_21.INJECT1_0 = "NO";
    defparam count_2674_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27027), .COUT(n27028), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_19.INJECT1_0 = "NO";
    defparam count_2674_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27026), .COUT(n27027), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_17.INJECT1_0 = "NO";
    defparam count_2674_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26641), .COUT(n26642));
    defparam sub_2068_add_2_15.INIT0 = 16'h5999;
    defparam sub_2068_add_2_15.INIT1 = 16'h5999;
    defparam sub_2068_add_2_15.INJECT1_0 = "NO";
    defparam sub_2068_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26640), .COUT(n26641));
    defparam sub_2068_add_2_13.INIT0 = 16'h5999;
    defparam sub_2068_add_2_13.INIT1 = 16'h5999;
    defparam sub_2068_add_2_13.INJECT1_0 = "NO";
    defparam sub_2068_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27025), .COUT(n27026), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_15.INJECT1_0 = "NO";
    defparam count_2674_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27024), .COUT(n27025), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_13.INJECT1_0 = "NO";
    defparam count_2674_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27023), .COUT(n27024), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_11.INJECT1_0 = "NO";
    defparam count_2674_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26639), .COUT(n26640));
    defparam sub_2068_add_2_11.INIT0 = 16'h5999;
    defparam sub_2068_add_2_11.INIT1 = 16'h5999;
    defparam sub_2068_add_2_11.INJECT1_0 = "NO";
    defparam sub_2068_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27022), .COUT(n27023), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_9.INJECT1_0 = "NO";
    defparam count_2674_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26638), .COUT(n26639));
    defparam sub_2068_add_2_9.INIT0 = 16'h5999;
    defparam sub_2068_add_2_9.INIT1 = 16'h5999;
    defparam sub_2068_add_2_9.INJECT1_0 = "NO";
    defparam sub_2068_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27021), .COUT(n27022), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_7.INJECT1_0 = "NO";
    defparam count_2674_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27020), .COUT(n27021), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_5.INJECT1_0 = "NO";
    defparam count_2674_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27019), .COUT(n27020), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_3.INJECT1_0 = "NO";
    defparam count_2674_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26637), .COUT(n26638));
    defparam sub_2068_add_2_7.INIT0 = 16'h5999;
    defparam sub_2068_add_2_7.INIT1 = 16'h5999;
    defparam sub_2068_add_2_7.INJECT1_0 = "NO";
    defparam sub_2068_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27019), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_1.INIT0 = 16'hF000;
    defparam count_2674_add_4_1.INIT1 = 16'h0555;
    defparam count_2674_add_4_1.INJECT1_0 = "NO";
    defparam count_2674_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26636), .COUT(n26637));
    defparam sub_2068_add_2_5.INIT0 = 16'h5999;
    defparam sub_2068_add_2_5.INIT1 = 16'h5999;
    defparam sub_2068_add_2_5.INJECT1_0 = "NO";
    defparam sub_2068_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26635), .COUT(n26636));
    defparam sub_2068_add_2_3.INIT0 = 16'h5999;
    defparam sub_2068_add_2_3.INIT1 = 16'h5999;
    defparam sub_2068_add_2_3.INJECT1_0 = "NO";
    defparam sub_2068_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2068_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26635));
    defparam sub_2068_add_2_1.INIT0 = 16'h0000;
    defparam sub_2068_add_2_1.INIT1 = 16'h5999;
    defparam sub_2068_add_2_1.INJECT1_0 = "NO";
    defparam sub_2068_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26634), .S1(n8159));
    defparam sub_2070_add_2_33.INIT0 = 16'h5999;
    defparam sub_2070_add_2_33.INIT1 = 16'h0000;
    defparam sub_2070_add_2_33.INJECT1_0 = "NO";
    defparam sub_2070_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26633), .COUT(n26634));
    defparam sub_2070_add_2_31.INIT0 = 16'h5999;
    defparam sub_2070_add_2_31.INIT1 = 16'h5999;
    defparam sub_2070_add_2_31.INJECT1_0 = "NO";
    defparam sub_2070_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26632), .COUT(n26633));
    defparam sub_2070_add_2_29.INIT0 = 16'h5999;
    defparam sub_2070_add_2_29.INIT1 = 16'h5999;
    defparam sub_2070_add_2_29.INJECT1_0 = "NO";
    defparam sub_2070_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26631), .COUT(n26632));
    defparam sub_2070_add_2_27.INIT0 = 16'h5999;
    defparam sub_2070_add_2_27.INIT1 = 16'h5999;
    defparam sub_2070_add_2_27.INJECT1_0 = "NO";
    defparam sub_2070_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26630), .COUT(n26631));
    defparam sub_2070_add_2_25.INIT0 = 16'h5999;
    defparam sub_2070_add_2_25.INIT1 = 16'h5999;
    defparam sub_2070_add_2_25.INJECT1_0 = "NO";
    defparam sub_2070_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26629), .COUT(n26630));
    defparam sub_2070_add_2_23.INIT0 = 16'h5999;
    defparam sub_2070_add_2_23.INIT1 = 16'h5999;
    defparam sub_2070_add_2_23.INJECT1_0 = "NO";
    defparam sub_2070_add_2_23.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (n2, databus, \read_value[10] , n8, n31425, \register_addr[0] , 
            read_value, read_value_adj_308, n46, n52, databus_out, 
            rw, read_value_adj_309, \read_value[10]_adj_157 , n52_adj_158, 
            n31446, n2_adj_159, \read_value[9]_adj_160 , n8_adj_161, 
            \read_value[9]_adj_162 , n2_adj_163, \select[7] , n176, 
            \read_value[8]_adj_164 , n8_adj_165, \register_addr[1] , n2_adj_166, 
            \read_value[24]_adj_167 , n8_adj_168, \read_value[24]_adj_169 , 
            \read_value[8]_adj_170 , n2_adj_171, \read_value[7]_adj_172 , 
            \read_value[7]_adj_173 , n31443, n3, read_value_adj_310, 
            n64, n66, read_value_adj_311, \read_value[14]_adj_190 , 
            n2_adj_191, \read_value[6]_adj_192 , \read_value[6]_adj_193 , 
            n3_adj_194, n2_adj_195, \read_value[5]_adj_196 , \read_value[5]_adj_197 , 
            n33384, n3_adj_198, n2_adj_199, \read_value[4]_adj_200 , 
            \read_value[4]_adj_201 , n3_adj_202, n2_adj_203, \read_value[3]_adj_204 , 
            \read_value[3]_adj_205 , n2_adj_206, \read_value[22]_adj_207 , 
            n8_adj_208, n3_adj_209, n2_adj_210, \read_value[2]_adj_211 , 
            \read_value[2]_adj_212 , \read_value[22]_adj_213 , n3_adj_214, 
            n10, \read_value[1]_adj_215 , n3_adj_216, \read_value[1]_adj_217 , 
            n2_adj_218, \read_value[13]_adj_219 , n8_adj_220, n2_adj_221, 
            \read_value[13]_adj_222 , \read_value[23]_adj_223 , n8_adj_224, 
            n2_adj_225, n2_adj_226, \read_value[12]_adj_227 , n8_adj_228, 
            \read_value[23]_adj_229 , \read_value[12]_adj_230 , \read_value[21]_adj_231 , 
            n8_adj_232, read_size, \select[1] , n13, n31482, n9, 
            \read_size[0]_adj_233 , n18, \read_size[0]_adj_234 , \read_size[0]_adj_235 , 
            n31464, \select[2] , n14, n31473, n5, \read_size[0]_adj_236 , 
            \read_size[0]_adj_237 , n31444, \select[5] , \read_size[0]_adj_238 , 
            n2_adj_239, \read_value[11]_adj_240 , n8_adj_241, n6, \read_size[2]_adj_242 , 
            \reg_size[2] , \read_size[2]_adj_243 , n9_adj_244, \read_size[2]_adj_245 , 
            n31470, \read_value[11]_adj_246 , \read_value[21]_adj_247 , 
            n2_adj_248, \read_value[25]_adj_249 , n8_adj_250, \read_value[25]_adj_251 , 
            \register_addr[2] , n2_adj_252, n2_adj_253, \read_value[20]_adj_254 , 
            n8_adj_255, \read_value[16]_adj_256 , n8_adj_257, n31587, 
            \sendcount[1] , n13155, n31456, \read_value[20]_adj_258 , 
            n2_adj_259, n2_adj_260, \read_value[0]_adj_261 , \read_value[0]_adj_262 , 
            n3_adj_263, n2_adj_264, \read_value[26]_adj_265 , n8_adj_266, 
            \read_value[26]_adj_267 , \read_value[16]_adj_268 , n2_adj_269, 
            \read_value[19]_adj_270 , n8_adj_271, n29236, n2_adj_272, 
            \read_value[19]_adj_273 , n2_adj_274, \read_value[18]_adj_275 , 
            n8_adj_276, n2_adj_277, \read_value[31]_adj_278 , n8_adj_279, 
            \read_value[14]_adj_280 , n8_adj_281, \read_value[31]_adj_282 , 
            n2_adj_283, \read_value[30]_adj_284 , n8_adj_285, \read_value[18]_adj_286 , 
            \read_value[30]_adj_287 , n2_adj_288, \read_value[17]_adj_289 , 
            \read_value[29]_adj_290 , n8_adj_291, \read_value[29]_adj_292 , 
            n2_adj_293, n2_adj_294, \read_value[15]_adj_295 , n8_adj_296, 
            \read_value[28]_adj_297 , n8_adj_298, \read_value[17]_adj_299 , 
            n8_adj_300, \read_value[28]_adj_301 , n2_adj_302, \read_value[27]_adj_303 , 
            n8_adj_304, \read_value[15]_adj_305 , \read_value[27]_adj_306 , 
            GND_net, debug_c_c, n33386, rc_ch8_c, n29817, n33385, 
            n13956, n27563, n29783, rc_ch7_c, n33387, n27542, n29826, 
            rc_ch4_c, n27549, n29837, rc_ch3_c, n14499, n27540, 
            n29839, n29529, n29943, n14_adj_307, n29831, rc_ch2_c, 
            n31411, n14512, n29846, n27535, n31511, n14513, rc_ch1_c, 
            n29829, n27546, n29810) /* synthesis syn_module_defined=1 */ ;
    input n2;
    output [31:0]databus;
    input \read_value[10] ;
    input n8;
    input n31425;
    input \register_addr[0] ;
    input [31:0]read_value;
    input [31:0]read_value_adj_308;
    input n46;
    input n52;
    input [31:0]databus_out;
    input rw;
    input [31:0]read_value_adj_309;
    input \read_value[10]_adj_157 ;
    input n52_adj_158;
    input n31446;
    input n2_adj_159;
    input \read_value[9]_adj_160 ;
    input n8_adj_161;
    input \read_value[9]_adj_162 ;
    input n2_adj_163;
    input \select[7] ;
    input n176;
    input \read_value[8]_adj_164 ;
    input n8_adj_165;
    input \register_addr[1] ;
    input n2_adj_166;
    input \read_value[24]_adj_167 ;
    input n8_adj_168;
    input \read_value[24]_adj_169 ;
    input \read_value[8]_adj_170 ;
    input n2_adj_171;
    input \read_value[7]_adj_172 ;
    input \read_value[7]_adj_173 ;
    input n31443;
    input n3;
    input [7:0]read_value_adj_310;
    input n64;
    input n66;
    input [7:0]read_value_adj_311;
    input \read_value[14]_adj_190 ;
    input n2_adj_191;
    input \read_value[6]_adj_192 ;
    input \read_value[6]_adj_193 ;
    input n3_adj_194;
    input n2_adj_195;
    input \read_value[5]_adj_196 ;
    input \read_value[5]_adj_197 ;
    input n33384;
    input n3_adj_198;
    input n2_adj_199;
    input \read_value[4]_adj_200 ;
    input \read_value[4]_adj_201 ;
    input n3_adj_202;
    input n2_adj_203;
    input \read_value[3]_adj_204 ;
    input \read_value[3]_adj_205 ;
    input n2_adj_206;
    input \read_value[22]_adj_207 ;
    input n8_adj_208;
    input n3_adj_209;
    input n2_adj_210;
    input \read_value[2]_adj_211 ;
    input \read_value[2]_adj_212 ;
    input \read_value[22]_adj_213 ;
    input n3_adj_214;
    input n10;
    input \read_value[1]_adj_215 ;
    input n3_adj_216;
    input \read_value[1]_adj_217 ;
    input n2_adj_218;
    input \read_value[13]_adj_219 ;
    input n8_adj_220;
    input n2_adj_221;
    input \read_value[13]_adj_222 ;
    input \read_value[23]_adj_223 ;
    input n8_adj_224;
    input n2_adj_225;
    input n2_adj_226;
    input \read_value[12]_adj_227 ;
    input n8_adj_228;
    input \read_value[23]_adj_229 ;
    input \read_value[12]_adj_230 ;
    input \read_value[21]_adj_231 ;
    input n8_adj_232;
    input [2:0]read_size;
    input \select[1] ;
    output n13;
    input n31482;
    input n9;
    input \read_size[0]_adj_233 ;
    output n18;
    input \read_size[0]_adj_234 ;
    input \read_size[0]_adj_235 ;
    input n31464;
    input \select[2] ;
    output n14;
    input n31473;
    input n5;
    input \read_size[0]_adj_236 ;
    input \read_size[0]_adj_237 ;
    input n31444;
    input \select[5] ;
    input \read_size[0]_adj_238 ;
    input n2_adj_239;
    input \read_value[11]_adj_240 ;
    input n8_adj_241;
    input n6;
    input \read_size[2]_adj_242 ;
    output \reg_size[2] ;
    input \read_size[2]_adj_243 ;
    input n9_adj_244;
    input \read_size[2]_adj_245 ;
    input n31470;
    input \read_value[11]_adj_246 ;
    input \read_value[21]_adj_247 ;
    input n2_adj_248;
    input \read_value[25]_adj_249 ;
    input n8_adj_250;
    input \read_value[25]_adj_251 ;
    input \register_addr[2] ;
    input n2_adj_252;
    input n2_adj_253;
    input \read_value[20]_adj_254 ;
    input n8_adj_255;
    input \read_value[16]_adj_256 ;
    input n8_adj_257;
    output n31587;
    input \sendcount[1] ;
    output n13155;
    input n31456;
    input \read_value[20]_adj_258 ;
    input n2_adj_259;
    input n2_adj_260;
    input \read_value[0]_adj_261 ;
    input \read_value[0]_adj_262 ;
    input n3_adj_263;
    input n2_adj_264;
    input \read_value[26]_adj_265 ;
    input n8_adj_266;
    input \read_value[26]_adj_267 ;
    input \read_value[16]_adj_268 ;
    input n2_adj_269;
    input \read_value[19]_adj_270 ;
    input n8_adj_271;
    output n29236;
    input n2_adj_272;
    input \read_value[19]_adj_273 ;
    input n2_adj_274;
    input \read_value[18]_adj_275 ;
    input n8_adj_276;
    input n2_adj_277;
    input \read_value[31]_adj_278 ;
    input n8_adj_279;
    input \read_value[14]_adj_280 ;
    input n8_adj_281;
    input \read_value[31]_adj_282 ;
    input n2_adj_283;
    input \read_value[30]_adj_284 ;
    input n8_adj_285;
    input \read_value[18]_adj_286 ;
    input \read_value[30]_adj_287 ;
    input n2_adj_288;
    input \read_value[17]_adj_289 ;
    input \read_value[29]_adj_290 ;
    input n8_adj_291;
    input \read_value[29]_adj_292 ;
    input n2_adj_293;
    input n2_adj_294;
    input \read_value[15]_adj_295 ;
    input n8_adj_296;
    input \read_value[28]_adj_297 ;
    input n8_adj_298;
    input \read_value[17]_adj_299 ;
    input n8_adj_300;
    input \read_value[28]_adj_301 ;
    input n2_adj_302;
    input \read_value[27]_adj_303 ;
    input n8_adj_304;
    input \read_value[15]_adj_305 ;
    input \read_value[27]_adj_306 ;
    input GND_net;
    input debug_c_c;
    input n33386;
    input rc_ch8_c;
    output n29817;
    input n33385;
    input n13956;
    input n27563;
    output n29783;
    input rc_ch7_c;
    input n33387;
    input n27542;
    output n29826;
    input rc_ch4_c;
    input n27549;
    output n29837;
    input rc_ch3_c;
    input n14499;
    input n27540;
    output n29839;
    output n29529;
    output n29943;
    input n14_adj_307;
    output n29831;
    input rc_ch2_c;
    input n31411;
    input n14512;
    output n29846;
    input n27535;
    input n31511;
    input n14513;
    input rc_ch1_c;
    output n29829;
    input n27546;
    output n29810;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n13_c, n11, n5_c, n10_c;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n30332, n13_adj_224, n11_adj_225, n5_adj_227, n10_adj_228, 
        n13_adj_234, n11_adj_235, n5_adj_237;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(211[12:21])
    
    wire n10_adj_238, n30777, n30776, n30778;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n30336, n13_adj_240, n11_adj_241, n5_adj_243, n10_adj_244;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n30779, n1209, n30780, n15, n20, n7;
    wire [7:0]read_value_adj_588;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(210[12:22])
    
    wire n18_c, n12, n46_adj_257, n14_c, n5_adj_263, n10_adj_265, 
        n30815, n15_adj_266, n20_adj_267, n7_adj_269, n30816, n18_adj_272, 
        n12_adj_273, n14_adj_275, n30818, n15_adj_281, n20_adj_282, 
        n7_adj_284, n18_adj_287, n12_adj_288, n14_adj_290, n1224, 
        n30819, n15_adj_296, n20_adj_297, n7_adj_299, n18_adj_302, 
        n12_adj_303, n31156, n31154, n1239, n31157, n31153, n14_adj_305, 
        n15_adj_311, n20_adj_312, n7_adj_314, n18_adj_317, n12_adj_318, 
        n13_adj_319, n11_adj_320, n5_adj_322, n10_adj_323, n14_adj_328, 
        n30837, n30838, n15_adj_334, n20_adj_335, n7_adj_337, n30840, 
        n18_adj_340, n12_adj_341, n14_adj_345, n1194, n30841, n19, 
        n8_adj_351, n18_adj_352, n12_adj_353, n16, n14_adj_356, n13_adj_364, 
        n11_adj_365, n5_adj_367, n10_adj_368, n13_adj_370, n11_adj_371, 
        n5_adj_373, n10_adj_378, n30333, n13_adj_382, n11_adj_383, 
        n5_adj_385, n13_adj_386, n11_adj_387, n5_adj_389, n10_adj_390, 
        n10_adj_398, n16_adj_402, n12_adj_408, n13_adj_415, n11_adj_416, 
        n5_adj_418, n10_adj_419, n10_adj_423, n8_adj_425, n30887, 
        n30884, n30885, n1179, n30888, n31304, n31303, n31306, 
        n31307, n13_adj_433, n11_adj_434, n5_adj_436, n31316, n10_adj_437, 
        n31315, n31320, n31317, n31321, n31318, n31319, n1164, 
        n13_adj_443, n11_adj_444, n5_adj_446, n13_adj_447, n11_adj_448, 
        n5_adj_450, n10_adj_451, n10_adj_453, n31308, n31305, n31309, 
        n30890, n30843, n30782, n30338, n30821, n31159, n13_adj_461, 
        n11_adj_462, n15_adj_464, n20_adj_465, n7_adj_467, n18_adj_470, 
        n12_adj_471, n14_adj_473, n13_adj_475, n11_adj_476, n5_adj_478, 
        n10_adj_481, n30337, n30334, n31158, n31155, n13_adj_491, 
        n11_adj_492, n5_adj_494, n10_adj_495, n30335, n13_adj_499, 
        n11_adj_500, n5_adj_502, n30889, n30886, n13_adj_505, n11_adj_506, 
        n5_adj_508, n10_adj_509, n13_adj_513, n11_adj_514, n5_adj_516, 
        n10_adj_517, n5_adj_521, n13_adj_526, n11_adj_527, n5_adj_529, 
        n10_adj_530, n30842, n30839, n13_adj_538, n11_adj_539, n5_adj_541, 
        n10_adj_543, n10_adj_544, n13_adj_550, n11_adj_551, n5_adj_553, 
        n13_adj_556, n11_adj_557, n10_adj_559, n30820, n30817, n10_adj_563, 
        n13_adj_571, n11_adj_572, n5_adj_574, n10_adj_575, n30781;
    
    LUT4 i7_4_lut (.A(n13_c), .B(n11), .C(n2), .D(n5_c), .Z(databus[10])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut (.A(\read_value[10] ), .B(n10_c), .C(n8), .D(n31425), 
         .Z(n13_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_22610 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n30332)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22610.init = 16'h2222;
    LUT4 i3_4_lut (.A(read_value[10]), .B(read_value_adj_308[10]), .C(n46), 
         .D(n52), .Z(n11)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 Select_4282_i5_2_lut (.A(databus_out[10]), .B(rw), .Z(n5_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4282_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut (.A(read_value_adj_309[10]), .B(\read_value[10]_adj_157 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 i7_4_lut_adj_341 (.A(n13_adj_224), .B(n11_adj_225), .C(n2_adj_159), 
         .D(n5_adj_227), .Z(databus[9])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_341.init = 16'hfffe;
    LUT4 i5_4_lut_adj_342 (.A(\read_value[9]_adj_160 ), .B(n10_adj_228), 
         .C(n8_adj_161), .D(n31425), .Z(n13_adj_224)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_342.init = 16'hfefc;
    LUT4 i3_4_lut_adj_343 (.A(read_value[9]), .B(read_value_adj_308[9]), 
         .C(n46), .D(n52), .Z(n11_adj_225)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_343.init = 16'heca0;
    LUT4 Select_4285_i5_2_lut (.A(databus_out[9]), .B(rw), .Z(n5_adj_227)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4285_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_344 (.A(read_value_adj_309[9]), .B(\read_value[9]_adj_162 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_228)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_344.init = 16'heca0;
    LUT4 i7_4_lut_adj_345 (.A(n13_adj_234), .B(n11_adj_235), .C(n2_adj_163), 
         .D(n5_adj_237), .Z(databus[8])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_345.init = 16'hfffe;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_346 (.A(\read_value[8]_adj_164 ), .B(n10_adj_238), 
         .C(n8_adj_165), .D(n31425), .Z(n13_adj_234)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_346.init = 16'hfefc;
    PFUMX i22677 (.BLUT(n30777), .ALUT(n30776), .C0(\register_addr[1] ), 
          .Z(n30778));
    LUT4 \register_1[[5__bdd_2_lut_22781  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n30336)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_22781 .init = 16'h8888;
    LUT4 i7_4_lut_adj_347 (.A(n13_adj_240), .B(n11_adj_241), .C(n2_adj_166), 
         .D(n5_adj_243), .Z(databus[24])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_347.init = 16'hfffe;
    LUT4 i5_4_lut_adj_348 (.A(\read_value[24]_adj_167 ), .B(n10_adj_244), 
         .C(n8_adj_168), .D(n31425), .Z(n13_adj_240)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_348.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_22695 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n30777)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22695.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_22694 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n30776)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22694.init = 16'h2222;
    LUT4 i3_4_lut_adj_349 (.A(read_value[24]), .B(read_value_adj_308[24]), 
         .C(n46), .D(n52), .Z(n11_adj_241)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_349.init = 16'heca0;
    LUT4 n1209_bdd_3_lut_22679 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n30779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1209_bdd_3_lut_22679.init = 16'hcaca;
    LUT4 Select_4240_i5_2_lut (.A(databus_out[24]), .B(rw), .Z(n5_adj_243)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4240_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_350 (.A(read_value_adj_309[24]), .B(\read_value[24]_adj_169 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_244)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_350.init = 16'heca0;
    LUT4 n1209_bdd_3_lut_22974 (.A(n1209), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n30780)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1209_bdd_3_lut_22974.init = 16'he2e2;
    LUT4 i3_4_lut_adj_351 (.A(read_value[8]), .B(read_value_adj_308[8]), 
         .C(n46), .D(n52), .Z(n11_adj_235)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_351.init = 16'heca0;
    LUT4 Select_4288_i5_2_lut (.A(databus_out[8]), .B(rw), .Z(n5_adj_237)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4288_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_352 (.A(read_value_adj_309[8]), .B(\read_value[8]_adj_170 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_238)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_352.init = 16'heca0;
    LUT4 i10_4_lut (.A(n15), .B(n20), .C(n2_adj_171), .D(n7), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i4_4_lut (.A(\read_value[7]_adj_172 ), .B(\read_value[7]_adj_173 ), 
         .C(n31446), .D(n31443), .Z(n15)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut.init = 16'heca0;
    LUT4 i9_4_lut (.A(read_value_adj_588[7]), .B(n18_c), .C(n12), .D(n46_adj_257), 
         .Z(n20)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut.init = 16'hfefc;
    LUT4 Select_4289_i7_2_lut (.A(databus_out[7]), .B(rw), .Z(n7)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4289_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_353 (.A(read_value[7]), .B(n14_c), .C(n3), .D(n46), 
         .Z(n18_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_353.init = 16'hfefc;
    LUT4 i1_4_lut (.A(read_value_adj_308[7]), .B(read_value_adj_310[7]), 
         .C(n52), .D(n64), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i3_4_lut_adj_354 (.A(read_value_adj_309[7]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[7]), .Z(n14_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_354.init = 16'heca0;
    LUT4 i14_2_lut (.A(\select[7] ), .B(rw), .Z(n46_adj_257)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam i14_2_lut.init = 16'h8888;
    LUT4 Select_4270_i5_2_lut (.A(databus_out[14]), .B(rw), .Z(n5_adj_263)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4270_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_355 (.A(read_value_adj_309[14]), .B(\read_value[14]_adj_190 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_265)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_355.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22705 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n30815)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22705.init = 16'h2222;
    LUT4 i10_4_lut_adj_356 (.A(n15_adj_266), .B(n20_adj_267), .C(n2_adj_191), 
         .D(n7_adj_269), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_356.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_22706 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n30816)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22706.init = 16'he4e4;
    LUT4 i4_4_lut_adj_357 (.A(\read_value[6]_adj_192 ), .B(\read_value[6]_adj_193 ), 
         .C(n31446), .D(n31443), .Z(n15_adj_266)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_357.init = 16'heca0;
    LUT4 i9_4_lut_adj_358 (.A(read_value_adj_588[6]), .B(n18_adj_272), .C(n12_adj_273), 
         .D(n46_adj_257), .Z(n20_adj_267)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_358.init = 16'hfefc;
    LUT4 Select_4290_i7_2_lut (.A(databus_out[6]), .B(rw), .Z(n7_adj_269)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4290_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_359 (.A(read_value[6]), .B(n14_adj_275), .C(n3_adj_194), 
         .D(n46), .Z(n18_adj_272)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_359.init = 16'hfefc;
    LUT4 i1_4_lut_adj_360 (.A(read_value_adj_308[6]), .B(read_value_adj_310[6]), 
         .C(n52), .D(n64), .Z(n12_adj_273)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_360.init = 16'heca0;
    LUT4 i3_4_lut_adj_361 (.A(read_value_adj_309[6]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[6]), .Z(n14_adj_275)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_361.init = 16'heca0;
    LUT4 n1224_bdd_3_lut_22700 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n30818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1224_bdd_3_lut_22700.init = 16'hcaca;
    LUT4 i10_4_lut_adj_362 (.A(n15_adj_281), .B(n20_adj_282), .C(n2_adj_195), 
         .D(n7_adj_284), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_362.init = 16'hfffe;
    LUT4 i4_4_lut_adj_363 (.A(\read_value[5]_adj_196 ), .B(\read_value[5]_adj_197 ), 
         .C(n31446), .D(n31443), .Z(n15_adj_281)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_363.init = 16'heca0;
    LUT4 i9_4_lut_adj_364 (.A(read_value_adj_588[5]), .B(n18_adj_287), .C(n12_adj_288), 
         .D(n46_adj_257), .Z(n20_adj_282)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_364.init = 16'hfefc;
    LUT4 Select_4291_i7_2_lut (.A(databus_out[5]), .B(n33384), .Z(n7_adj_284)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4291_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_365 (.A(read_value[5]), .B(n14_adj_290), .C(n3_adj_198), 
         .D(n46), .Z(n18_adj_287)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_365.init = 16'hfefc;
    LUT4 i1_4_lut_adj_366 (.A(read_value_adj_308[5]), .B(read_value_adj_310[5]), 
         .C(n52), .D(n64), .Z(n12_adj_288)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_366.init = 16'heca0;
    LUT4 i3_4_lut_adj_367 (.A(read_value_adj_309[5]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[5]), .Z(n14_adj_290)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_367.init = 16'heca0;
    LUT4 n1224_bdd_3_lut_22963 (.A(n1224), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n30819)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1224_bdd_3_lut_22963.init = 16'he2e2;
    LUT4 i10_4_lut_adj_368 (.A(n15_adj_296), .B(n20_adj_297), .C(n2_adj_199), 
         .D(n7_adj_299), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_368.init = 16'hfffe;
    LUT4 i4_4_lut_adj_369 (.A(\read_value[4]_adj_200 ), .B(\read_value[4]_adj_201 ), 
         .C(n31446), .D(n31443), .Z(n15_adj_296)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_369.init = 16'heca0;
    LUT4 i9_4_lut_adj_370 (.A(read_value_adj_588[4]), .B(n18_adj_302), .C(n12_adj_303), 
         .D(n46_adj_257), .Z(n20_adj_297)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_370.init = 16'hfefc;
    LUT4 n1239_bdd_3_lut_22871 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n31156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1239_bdd_3_lut_22871.init = 16'hcaca;
    LUT4 Select_4292_i7_2_lut (.A(databus_out[4]), .B(n33384), .Z(n7_adj_299)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4292_i7_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_22929 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n31154)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22929.init = 16'he4e4;
    LUT4 n1239_bdd_3_lut_23345 (.A(n1239), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n31157)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1239_bdd_3_lut_23345.init = 16'he2e2;
    LUT4 register_addr_1__bdd_2_lut_22928 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n31153)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22928.init = 16'h2222;
    LUT4 i7_4_lut_adj_371 (.A(read_value[4]), .B(n14_adj_305), .C(n3_adj_202), 
         .D(n46), .Z(n18_adj_302)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_371.init = 16'hfefc;
    LUT4 i1_4_lut_adj_372 (.A(read_value_adj_308[4]), .B(read_value_adj_310[4]), 
         .C(n52), .D(n64), .Z(n12_adj_303)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_372.init = 16'heca0;
    LUT4 i3_4_lut_adj_373 (.A(read_value_adj_309[4]), .B(read_value_adj_311[4]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_305)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_373.init = 16'heca0;
    LUT4 i10_4_lut_adj_374 (.A(n15_adj_311), .B(n20_adj_312), .C(n2_adj_203), 
         .D(n7_adj_314), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_374.init = 16'hfffe;
    LUT4 i4_4_lut_adj_375 (.A(\read_value[3]_adj_204 ), .B(\read_value[3]_adj_205 ), 
         .C(n31446), .D(n31443), .Z(n15_adj_311)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_375.init = 16'heca0;
    LUT4 i9_4_lut_adj_376 (.A(read_value_adj_588[3]), .B(n18_adj_317), .C(n12_adj_318), 
         .D(n46_adj_257), .Z(n20_adj_312)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_376.init = 16'hfefc;
    LUT4 i7_4_lut_adj_377 (.A(n13_adj_319), .B(n11_adj_320), .C(n2_adj_206), 
         .D(n5_adj_322), .Z(databus[22])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_377.init = 16'hfffe;
    LUT4 i5_4_lut_adj_378 (.A(\read_value[22]_adj_207 ), .B(n10_adj_323), 
         .C(n8_adj_208), .D(n31425), .Z(n13_adj_319)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_378.init = 16'hfefc;
    LUT4 i3_4_lut_adj_379 (.A(read_value[22]), .B(read_value_adj_308[22]), 
         .C(n46), .D(n52), .Z(n11_adj_320)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_379.init = 16'heca0;
    LUT4 Select_4293_i7_2_lut (.A(databus_out[3]), .B(n33384), .Z(n7_adj_314)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4293_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_380 (.A(read_value[3]), .B(n14_adj_328), .C(n3_adj_209), 
         .D(n46), .Z(n18_adj_317)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_380.init = 16'hfefc;
    LUT4 i1_4_lut_adj_381 (.A(read_value_adj_308[3]), .B(read_value_adj_310[3]), 
         .C(n52), .D(n64), .Z(n12_adj_318)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_381.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22742 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n30837)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22742.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_22743 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n30838)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22743.init = 16'he4e4;
    LUT4 i3_4_lut_adj_382 (.A(read_value_adj_309[3]), .B(read_value_adj_311[3]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_328)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_382.init = 16'heca0;
    LUT4 i10_4_lut_adj_383 (.A(n15_adj_334), .B(n20_adj_335), .C(n2_adj_210), 
         .D(n7_adj_337), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_383.init = 16'hfffe;
    LUT4 n1194_bdd_3_lut_22715 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n30840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1194_bdd_3_lut_22715.init = 16'hcaca;
    LUT4 Select_4246_i5_2_lut (.A(databus_out[22]), .B(rw), .Z(n5_adj_322)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4246_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_384 (.A(\read_value[2]_adj_211 ), .B(\read_value[2]_adj_212 ), 
         .C(n31446), .D(n31443), .Z(n15_adj_334)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_384.init = 16'heca0;
    LUT4 i9_4_lut_adj_385 (.A(read_value_adj_588[2]), .B(n18_adj_340), .C(n12_adj_341), 
         .D(n46_adj_257), .Z(n20_adj_335)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_385.init = 16'hfefc;
    LUT4 Select_4294_i7_2_lut (.A(databus_out[2]), .B(n33384), .Z(n7_adj_337)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4294_i7_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_386 (.A(read_value_adj_309[22]), .B(\read_value[22]_adj_213 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_323)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_386.init = 16'heca0;
    LUT4 i7_4_lut_adj_387 (.A(read_value[2]), .B(n14_adj_345), .C(n3_adj_214), 
         .D(n46), .Z(n18_adj_340)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_387.init = 16'hfefc;
    LUT4 i1_4_lut_adj_388 (.A(read_value_adj_308[2]), .B(read_value_adj_310[2]), 
         .C(n52), .D(n64), .Z(n12_adj_341)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_388.init = 16'heca0;
    LUT4 i3_4_lut_adj_389 (.A(read_value_adj_309[2]), .B(read_value_adj_311[2]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_345)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_389.init = 16'heca0;
    LUT4 n1194_bdd_3_lut_22940 (.A(n1194), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n30841)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1194_bdd_3_lut_22940.init = 16'he2e2;
    LUT4 i10_4_lut_adj_390 (.A(n19), .B(n8_adj_351), .C(n18_adj_352), 
         .D(n12_adj_353), .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_390.init = 16'hfffe;
    LUT4 i8_4_lut (.A(read_value_adj_588[1]), .B(n16), .C(n10), .D(n46_adj_257), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut.init = 16'hfefc;
    LUT4 Select_4295_i8_2_lut (.A(databus_out[1]), .B(rw), .Z(n8_adj_351)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4295_i8_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_391 (.A(\read_value[1]_adj_215 ), .B(n14_adj_356), 
         .C(n3_adj_216), .D(n31443), .Z(n18_adj_352)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_391.init = 16'hfefc;
    LUT4 i1_4_lut_adj_392 (.A(read_value_adj_308[1]), .B(read_value_adj_310[1]), 
         .C(n52), .D(n64), .Z(n12_adj_353)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_392.init = 16'heca0;
    LUT4 i5_4_lut_adj_393 (.A(\read_value[1]_adj_217 ), .B(read_value[1]), 
         .C(n31425), .D(n46), .Z(n16)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i5_4_lut_adj_393.init = 16'heca0;
    LUT4 i3_4_lut_adj_394 (.A(read_value_adj_309[1]), .B(read_value_adj_311[1]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_356)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_394.init = 16'heca0;
    LUT4 i7_4_lut_adj_395 (.A(n13_adj_364), .B(n11_adj_365), .C(n2_adj_218), 
         .D(n5_adj_367), .Z(databus[13])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_395.init = 16'hfffe;
    LUT4 i5_4_lut_adj_396 (.A(\read_value[13]_adj_219 ), .B(n10_adj_368), 
         .C(n8_adj_220), .D(n31425), .Z(n13_adj_364)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_396.init = 16'hfefc;
    LUT4 i7_4_lut_adj_397 (.A(n13_adj_370), .B(n11_adj_371), .C(n2_adj_221), 
         .D(n5_adj_373), .Z(databus[23])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_397.init = 16'hfffe;
    LUT4 i3_4_lut_adj_398 (.A(read_value[13]), .B(read_value_adj_308[13]), 
         .C(n46), .D(n52), .Z(n11_adj_365)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_398.init = 16'heca0;
    LUT4 Select_4273_i5_2_lut (.A(databus_out[13]), .B(n33384), .Z(n5_adj_367)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4273_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_399 (.A(read_value_adj_309[13]), .B(\read_value[13]_adj_222 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_368)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_399.init = 16'heca0;
    LUT4 i5_4_lut_adj_400 (.A(\read_value[23]_adj_223 ), .B(n10_adj_378), 
         .C(n8_adj_224), .D(n31425), .Z(n13_adj_370)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_400.init = 16'hfefc;
    LUT4 i3_4_lut_adj_401 (.A(read_value[23]), .B(read_value_adj_308[23]), 
         .C(n46), .D(n52), .Z(n11_adj_371)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_401.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_22584 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n30333)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22584.init = 16'he4e4;
    LUT4 i7_4_lut_adj_402 (.A(n13_adj_382), .B(n11_adj_383), .C(n2_adj_225), 
         .D(n5_adj_385), .Z(databus[21])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_402.init = 16'hfffe;
    LUT4 Select_4243_i5_2_lut (.A(databus_out[23]), .B(rw), .Z(n5_adj_373)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4243_i5_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_403 (.A(n13_adj_386), .B(n11_adj_387), .C(n2_adj_226), 
         .D(n5_adj_389), .Z(databus[12])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_403.init = 16'hfffe;
    LUT4 i5_4_lut_adj_404 (.A(\read_value[12]_adj_227 ), .B(n10_adj_390), 
         .C(n8_adj_228), .D(n31425), .Z(n13_adj_386)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_404.init = 16'hfefc;
    LUT4 i2_4_lut_adj_405 (.A(read_value_adj_309[23]), .B(\read_value[23]_adj_229 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_378)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_405.init = 16'heca0;
    LUT4 i3_4_lut_adj_406 (.A(read_value[12]), .B(read_value_adj_308[12]), 
         .C(n46), .D(n52), .Z(n11_adj_387)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_406.init = 16'heca0;
    LUT4 Select_4276_i5_2_lut (.A(databus_out[12]), .B(n33384), .Z(n5_adj_389)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4276_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_407 (.A(read_value_adj_309[12]), .B(\read_value[12]_adj_230 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_390)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_407.init = 16'heca0;
    LUT4 i5_4_lut_adj_408 (.A(\read_value[21]_adj_231 ), .B(n10_adj_398), 
         .C(n8_adj_232), .D(n31425), .Z(n13_adj_382)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_408.init = 16'hfefc;
    LUT4 i3_4_lut_adj_409 (.A(read_size[0]), .B(read_size_c[0]), .C(\select[1] ), 
         .D(\select[7] ), .Z(n13)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_409.init = 16'heca0;
    LUT4 i8_4_lut_adj_410 (.A(n31482), .B(n16_adj_402), .C(n9), .D(\read_size[0]_adj_233 ), 
         .Z(n18)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_410.init = 16'hfefc;
    LUT4 i4_4_lut_adj_411 (.A(\read_size[0]_adj_234 ), .B(\read_size[0]_adj_235 ), 
         .C(n31464), .D(\select[2] ), .Z(n14)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_411.init = 16'heca0;
    LUT4 i6_4_lut (.A(n31473), .B(n12_adj_408), .C(n5), .D(\read_size[0]_adj_236 ), 
         .Z(n16_adj_402)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 i3_4_lut_adj_412 (.A(read_value[21]), .B(read_value_adj_308[21]), 
         .C(n46), .D(n52), .Z(n11_adj_383)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_412.init = 16'heca0;
    LUT4 i2_4_lut_adj_413 (.A(\read_size[0]_adj_237 ), .B(n31444), .C(\select[5] ), 
         .D(\read_size[0]_adj_238 ), .Z(n12_adj_408)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_413.init = 16'heca0;
    LUT4 i7_4_lut_adj_414 (.A(n13_adj_415), .B(n11_adj_416), .C(n2_adj_239), 
         .D(n5_adj_418), .Z(databus[11])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_414.init = 16'hfffe;
    LUT4 i5_4_lut_adj_415 (.A(\read_value[11]_adj_240 ), .B(n10_adj_419), 
         .C(n8_adj_241), .D(n31425), .Z(n13_adj_415)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_415.init = 16'hfefc;
    LUT4 i3_4_lut_adj_416 (.A(read_value[11]), .B(read_value_adj_308[11]), 
         .C(n46), .D(n52), .Z(n11_adj_416)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_416.init = 16'heca0;
    LUT4 i5_4_lut_adj_417 (.A(n31444), .B(n10_adj_423), .C(n6), .D(\read_size[2]_adj_242 ), 
         .Z(\reg_size[2] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_417.init = 16'hfefc;
    LUT4 i4_4_lut_adj_418 (.A(\read_size[2]_adj_243 ), .B(n8_adj_425), .C(n9_adj_244), 
         .D(n31482), .Z(n10_adj_423)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_418.init = 16'hfefc;
    LUT4 n1179_bdd_3_lut_22748 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n30887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1179_bdd_3_lut_22748.init = 16'hcaca;
    LUT4 i2_4_lut_adj_419 (.A(read_size[2]), .B(\read_size[2]_adj_245 ), 
         .C(\select[1] ), .D(n31470), .Z(n8_adj_425)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_419.init = 16'heca0;
    LUT4 Select_4279_i5_2_lut (.A(databus_out[11]), .B(n33384), .Z(n5_adj_418)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4279_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_420 (.A(read_value_adj_309[11]), .B(\read_value[11]_adj_246 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_419)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_420.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22787 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n30884)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22787.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_22788 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n30885)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22788.init = 16'he4e4;
    LUT4 n1179_bdd_3_lut_22912 (.A(n1179), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n30888)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1179_bdd_3_lut_22912.init = 16'he2e2;
    LUT4 Select_4249_i5_2_lut (.A(databus_out[21]), .B(rw), .Z(n5_adj_385)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4249_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_421 (.A(read_value_adj_309[21]), .B(\read_value[21]_adj_247 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_398)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_421.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_22951 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n31304)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22951.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_22950 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n31303)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22950.init = 16'h2222;
    LUT4 \register_1[[4__bdd_3_lut_23197  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n31306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_23197 .init = 16'hcaca;
    LUT4 \register_1[[4__bdd_2_lut_23198  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n31307)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_23198 .init = 16'h8888;
    LUT4 i7_4_lut_adj_422 (.A(n13_adj_433), .B(n11_adj_434), .C(n2_adj_248), 
         .D(n5_adj_436), .Z(databus[25])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_422.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n31316)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    LUT4 i5_4_lut_adj_423 (.A(\read_value[25]_adj_249 ), .B(n10_adj_437), 
         .C(n8_adj_250), .D(n31425), .Z(n13_adj_433)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_423.init = 16'hfefc;
    LUT4 i3_4_lut_adj_424 (.A(read_value[25]), .B(read_value_adj_308[25]), 
         .C(n46), .D(n52), .Z(n11_adj_434)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_424.init = 16'heca0;
    LUT4 Select_4237_i5_2_lut (.A(databus_out[25]), .B(rw), .Z(n5_adj_436)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4237_i5_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n31315)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_425 (.A(read_value_adj_309[25]), .B(\read_value[25]_adj_251 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_437)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_425.init = 16'heca0;
    L6MUX21 i22957 (.D0(n31320), .D1(n31317), .SD(\register_addr[2] ), 
            .Z(n31321));
    LUT4 n1164_bdd_3_lut_22954 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n31318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1164_bdd_3_lut_22954.init = 16'hcaca;
    PFUMX i22955 (.BLUT(n31319), .ALUT(n31318), .C0(\register_addr[1] ), 
          .Z(n31320));
    LUT4 n1164_bdd_3_lut_23161 (.A(n1164), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n31319)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1164_bdd_3_lut_23161.init = 16'he2e2;
    LUT4 i7_4_lut_adj_426 (.A(n13_adj_443), .B(n11_adj_444), .C(n2_adj_252), 
         .D(n5_adj_446), .Z(databus[20])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_426.init = 16'hfffe;
    PFUMX i22952 (.BLUT(n31316), .ALUT(n31315), .C0(\register_addr[1] ), 
          .Z(n31317));
    LUT4 i7_4_lut_adj_427 (.A(n13_adj_447), .B(n11_adj_448), .C(n2_adj_253), 
         .D(n5_adj_450), .Z(databus[16])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_427.init = 16'hfffe;
    LUT4 i5_4_lut_adj_428 (.A(\read_value[20]_adj_254 ), .B(n10_adj_451), 
         .C(n8_adj_255), .D(n31425), .Z(n13_adj_443)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_428.init = 16'hfefc;
    LUT4 i5_4_lut_adj_429 (.A(\read_value[16]_adj_256 ), .B(n10_adj_453), 
         .C(n8_adj_257), .D(n31425), .Z(n13_adj_447)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_429.init = 16'hfefc;
    L6MUX21 i22948 (.D0(n31308), .D1(n31305), .SD(\register_addr[2] ), 
            .Z(n31309));
    PFUMX i22946 (.BLUT(n31307), .ALUT(n31306), .C0(\register_addr[1] ), 
          .Z(n31308));
    LUT4 i3_4_lut_adj_430 (.A(read_value[20]), .B(read_value_adj_308[20]), 
         .C(n46), .D(n52), .Z(n11_adj_444)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_430.init = 16'heca0;
    LUT4 Select_4306_i1_2_lut_rep_444 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n31587)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4306_i1_2_lut_rep_444.init = 16'h8888;
    LUT4 i3_4_lut_adj_431 (.A(read_value[16]), .B(read_value_adj_308[16]), 
         .C(n46), .D(n52), .Z(n11_adj_448)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_431.init = 16'heca0;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n13155)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 Select_4264_i5_2_lut (.A(databus_out[16]), .B(n33384), .Z(n5_adj_450)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4264_i5_2_lut.init = 16'h2222;
    FD1S3IX read_value__i1 (.D(n30890), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n30843), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n30782), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n31309), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n30338), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(n30821), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i7 (.D(n31159), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i7.GSR = "ENABLED";
    PFUMX i22944 (.BLUT(n31304), .ALUT(n31303), .C0(\register_addr[1] ), 
          .Z(n31305));
    LUT4 Select_4252_i5_2_lut (.A(databus_out[20]), .B(rw), .Z(n5_adj_446)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4252_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_432 (.A(read_value_adj_309[20]), .B(\read_value[20]_adj_258 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_451)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_432.init = 16'heca0;
    LUT4 i7_4_lut_adj_433 (.A(n13_adj_461), .B(n11_adj_462), .C(n2_adj_259), 
         .D(n5_adj_263), .Z(databus[14])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_433.init = 16'hfffe;
    LUT4 i10_4_lut_adj_434 (.A(n15_adj_464), .B(n20_adj_465), .C(n2_adj_260), 
         .D(n7_adj_467), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_434.init = 16'hfffe;
    LUT4 i4_4_lut_adj_435 (.A(\read_value[0]_adj_261 ), .B(\read_value[0]_adj_262 ), 
         .C(n31446), .D(n31443), .Z(n15_adj_464)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_435.init = 16'heca0;
    LUT4 i9_4_lut_adj_436 (.A(read_value_adj_588[0]), .B(n18_adj_470), .C(n12_adj_471), 
         .D(n46_adj_257), .Z(n20_adj_465)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_436.init = 16'hfefc;
    LUT4 Select_4296_i7_2_lut (.A(databus_out[0]), .B(rw), .Z(n7_adj_467)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4296_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_437 (.A(read_value[0]), .B(n14_adj_473), .C(n3_adj_263), 
         .D(n46), .Z(n18_adj_470)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_437.init = 16'hfefc;
    LUT4 i7_4_lut_adj_438 (.A(n13_adj_475), .B(n11_adj_476), .C(n2_adj_264), 
         .D(n5_adj_478), .Z(databus[26])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_438.init = 16'hfffe;
    LUT4 i1_4_lut_adj_439 (.A(read_value_adj_308[0]), .B(read_value_adj_310[0]), 
         .C(n52), .D(n64), .Z(n12_adj_471)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_439.init = 16'heca0;
    LUT4 i5_4_lut_adj_440 (.A(\read_value[26]_adj_265 ), .B(n10_adj_481), 
         .C(n8_adj_266), .D(n31425), .Z(n13_adj_475)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_440.init = 16'hfefc;
    LUT4 i3_4_lut_adj_441 (.A(read_value_adj_309[0]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[0]), .Z(n14_adj_473)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_441.init = 16'heca0;
    LUT4 i3_4_lut_adj_442 (.A(read_value[26]), .B(read_value_adj_308[26]), 
         .C(n46), .D(n52), .Z(n11_adj_476)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_442.init = 16'heca0;
    LUT4 Select_4234_i5_2_lut (.A(databus_out[26]), .B(rw), .Z(n5_adj_478)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4234_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_443 (.A(read_value_adj_309[26]), .B(\read_value[26]_adj_267 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_481)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_443.init = 16'heca0;
    LUT4 i2_4_lut_adj_444 (.A(read_value_adj_309[16]), .B(\read_value[16]_adj_268 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_453)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_444.init = 16'heca0;
    L6MUX21 i22582 (.D0(n30337), .D1(n30334), .SD(\register_addr[2] ), 
            .Z(n30338));
    L6MUX21 i22874 (.D0(n31158), .D1(n31155), .SD(\register_addr[2] ), 
            .Z(n31159));
    PFUMX i22872 (.BLUT(n31157), .ALUT(n31156), .C0(\register_addr[1] ), 
          .Z(n31158));
    LUT4 i7_4_lut_adj_445 (.A(n13_adj_491), .B(n11_adj_492), .C(n2_adj_269), 
         .D(n5_adj_494), .Z(databus[19])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_445.init = 16'hfffe;
    PFUMX i22869 (.BLUT(n31154), .ALUT(n31153), .C0(\register_addr[1] ), 
          .Z(n31155));
    LUT4 i5_4_lut_adj_446 (.A(\read_value[19]_adj_270 ), .B(n10_adj_495), 
         .C(n8_adj_271), .D(n31425), .Z(n13_adj_491)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_446.init = 16'hfefc;
    LUT4 i1_2_lut (.A(\register_addr[0] ), .B(\register_addr[1] ), .Z(n29236)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    PFUMX i22580 (.BLUT(n30336), .ALUT(n30335), .C0(\register_addr[1] ), 
          .Z(n30337));
    LUT4 i3_4_lut_adj_447 (.A(read_value[19]), .B(read_value_adj_308[19]), 
         .C(n46), .D(n52), .Z(n11_adj_492)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_447.init = 16'heca0;
    FD1S3IX read_value__i0 (.D(n31321), .CK(\select[7] ), .CD(n31456), 
            .Q(read_value_adj_588[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=706, LSE_RLINE=718 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i7_4_lut_adj_448 (.A(n13_adj_499), .B(n11_adj_500), .C(n2_adj_272), 
         .D(n5_adj_502), .Z(databus[15])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_448.init = 16'hfffe;
    LUT4 Select_4255_i5_2_lut (.A(databus_out[19]), .B(rw), .Z(n5_adj_494)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4255_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_449 (.A(read_value_adj_309[19]), .B(\read_value[19]_adj_273 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_495)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_449.init = 16'heca0;
    L6MUX21 i22751 (.D0(n30889), .D1(n30886), .SD(\register_addr[2] ), 
            .Z(n30890));
    PFUMX i22749 (.BLUT(n30888), .ALUT(n30887), .C0(\register_addr[1] ), 
          .Z(n30889));
    LUT4 i7_4_lut_adj_450 (.A(n13_adj_505), .B(n11_adj_506), .C(n2_adj_274), 
         .D(n5_adj_508), .Z(databus[18])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_450.init = 16'hfffe;
    LUT4 i5_4_lut_adj_451 (.A(\read_value[18]_adj_275 ), .B(n10_adj_509), 
         .C(n8_adj_276), .D(n31425), .Z(n13_adj_505)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_451.init = 16'hfefc;
    LUT4 i3_4_lut_adj_452 (.A(read_value[18]), .B(read_value_adj_308[18]), 
         .C(n46), .D(n52), .Z(n11_adj_506)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_452.init = 16'heca0;
    PFUMX i22746 (.BLUT(n30885), .ALUT(n30884), .C0(\register_addr[1] ), 
          .Z(n30886));
    LUT4 i7_4_lut_adj_453 (.A(n13_adj_513), .B(n11_adj_514), .C(n2_adj_277), 
         .D(n5_adj_516), .Z(databus[31])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_453.init = 16'hfffe;
    LUT4 i5_4_lut_adj_454 (.A(\read_value[31]_adj_278 ), .B(n10_adj_517), 
         .C(n8_adj_279), .D(n31425), .Z(n13_adj_513)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_454.init = 16'hfefc;
    LUT4 i3_4_lut_adj_455 (.A(read_value[31]), .B(read_value_adj_308[31]), 
         .C(n46), .D(n52), .Z(n11_adj_514)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_455.init = 16'heca0;
    LUT4 Select_4261_i5_2_lut (.A(databus_out[17]), .B(n33384), .Z(n5_adj_521)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4261_i5_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_456 (.A(\read_value[14]_adj_280 ), .B(n10_adj_265), 
         .C(n8_adj_281), .D(n31425), .Z(n13_adj_461)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_456.init = 16'hfefc;
    LUT4 Select_4258_i5_2_lut (.A(databus_out[18]), .B(n33384), .Z(n5_adj_508)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4258_i5_2_lut.init = 16'h2222;
    LUT4 Select_4219_i5_2_lut (.A(databus_out[31]), .B(rw), .Z(n5_adj_516)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4219_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_457 (.A(read_value_adj_309[31]), .B(\read_value[31]_adj_282 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_517)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_457.init = 16'heca0;
    LUT4 i7_4_lut_adj_458 (.A(n13_adj_526), .B(n11_adj_527), .C(n2_adj_283), 
         .D(n5_adj_529), .Z(databus[30])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_458.init = 16'hfffe;
    LUT4 i5_4_lut_adj_459 (.A(\read_value[30]_adj_284 ), .B(n10_adj_530), 
         .C(n8_adj_285), .D(n31425), .Z(n13_adj_526)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_459.init = 16'hfefc;
    L6MUX21 i22718 (.D0(n30842), .D1(n30839), .SD(\register_addr[2] ), 
            .Z(n30843));
    LUT4 i3_4_lut_adj_460 (.A(read_value[30]), .B(read_value_adj_308[30]), 
         .C(n46), .D(n52), .Z(n11_adj_527)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_460.init = 16'heca0;
    LUT4 i2_4_lut_adj_461 (.A(read_value_adj_309[18]), .B(\read_value[18]_adj_286 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_509)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_461.init = 16'heca0;
    LUT4 Select_4222_i5_2_lut (.A(databus_out[30]), .B(rw), .Z(n5_adj_529)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4222_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_462 (.A(read_value_adj_309[30]), .B(\read_value[30]_adj_287 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_530)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_462.init = 16'heca0;
    PFUMX i22716 (.BLUT(n30841), .ALUT(n30840), .C0(\register_addr[1] ), 
          .Z(n30842));
    LUT4 \register_1[[5__bdd_3_lut_22780  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n30335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_22780 .init = 16'hcaca;
    LUT4 i7_4_lut_adj_463 (.A(n13_adj_538), .B(n11_adj_539), .C(n2_adj_288), 
         .D(n5_adj_541), .Z(databus[29])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_463.init = 16'hfffe;
    LUT4 i2_4_lut_adj_464 (.A(read_value_adj_309[17]), .B(\read_value[17]_adj_289 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_543)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_464.init = 16'heca0;
    LUT4 i5_4_lut_adj_465 (.A(\read_value[29]_adj_290 ), .B(n10_adj_544), 
         .C(n8_adj_291), .D(n31425), .Z(n13_adj_538)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_465.init = 16'hfefc;
    LUT4 i3_4_lut_adj_466 (.A(read_value[29]), .B(read_value_adj_308[29]), 
         .C(n46), .D(n52), .Z(n11_adj_539)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_466.init = 16'heca0;
    LUT4 Select_4225_i5_2_lut (.A(databus_out[29]), .B(rw), .Z(n5_adj_541)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4225_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_467 (.A(read_value_adj_309[29]), .B(\read_value[29]_adj_292 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_544)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_467.init = 16'heca0;
    PFUMX i22713 (.BLUT(n30838), .ALUT(n30837), .C0(\register_addr[1] ), 
          .Z(n30839));
    LUT4 i7_4_lut_adj_468 (.A(n13_adj_550), .B(n11_adj_551), .C(n2_adj_293), 
         .D(n5_adj_553), .Z(databus[28])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_468.init = 16'hfffe;
    LUT4 i3_4_lut_adj_469 (.A(read_value[14]), .B(read_value_adj_308[14]), 
         .C(n46), .D(n52), .Z(n11_adj_462)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_469.init = 16'heca0;
    LUT4 i7_4_lut_adj_470 (.A(n13_adj_556), .B(n11_adj_557), .C(n2_adj_294), 
         .D(n5_adj_521), .Z(databus[17])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_470.init = 16'hfffe;
    LUT4 i5_4_lut_adj_471 (.A(\read_value[15]_adj_295 ), .B(n10_adj_559), 
         .C(n8_adj_296), .D(n31425), .Z(n13_adj_499)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_471.init = 16'hfefc;
    L6MUX21 i22703 (.D0(n30820), .D1(n30817), .SD(\register_addr[2] ), 
            .Z(n30821));
    LUT4 i3_4_lut_adj_472 (.A(read_value[15]), .B(read_value_adj_308[15]), 
         .C(n46), .D(n52), .Z(n11_adj_500)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_472.init = 16'heca0;
    PFUMX i22701 (.BLUT(n30819), .ALUT(n30818), .C0(\register_addr[1] ), 
          .Z(n30820));
    PFUMX i22698 (.BLUT(n30816), .ALUT(n30815), .C0(\register_addr[1] ), 
          .Z(n30817));
    LUT4 i5_4_lut_adj_473 (.A(\read_value[28]_adj_297 ), .B(n10_adj_563), 
         .C(n8_adj_298), .D(n31425), .Z(n13_adj_550)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_473.init = 16'hfefc;
    LUT4 i3_4_lut_adj_474 (.A(read_value[28]), .B(read_value_adj_308[28]), 
         .C(n46), .D(n52), .Z(n11_adj_551)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_474.init = 16'heca0;
    LUT4 Select_4228_i5_2_lut (.A(databus_out[28]), .B(rw), .Z(n5_adj_553)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4228_i5_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_475 (.A(\read_value[17]_adj_299 ), .B(n10_adj_543), 
         .C(n8_adj_300), .D(n31425), .Z(n13_adj_556)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_475.init = 16'hfefc;
    LUT4 i2_4_lut_adj_476 (.A(read_value_adj_309[28]), .B(\read_value[28]_adj_301 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_563)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_476.init = 16'heca0;
    PFUMX i22578 (.BLUT(n30333), .ALUT(n30332), .C0(\register_addr[1] ), 
          .Z(n30334));
    LUT4 i7_4_lut_adj_477 (.A(n13_adj_571), .B(n11_adj_572), .C(n2_adj_302), 
         .D(n5_adj_574), .Z(databus[27])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_477.init = 16'hfffe;
    LUT4 i5_4_lut_adj_478 (.A(\read_value[27]_adj_303 ), .B(n10_adj_575), 
         .C(n8_adj_304), .D(n31425), .Z(n13_adj_571)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_478.init = 16'hfefc;
    LUT4 i3_4_lut_adj_479 (.A(read_value[27]), .B(read_value_adj_308[27]), 
         .C(n46), .D(n52), .Z(n11_adj_572)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_479.init = 16'heca0;
    L6MUX21 i22682 (.D0(n30781), .D1(n30778), .SD(\register_addr[2] ), 
            .Z(n30782));
    LUT4 i3_4_lut_adj_480 (.A(read_value[17]), .B(read_value_adj_308[17]), 
         .C(n46), .D(n52), .Z(n11_adj_557)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_480.init = 16'heca0;
    LUT4 Select_4267_i5_2_lut (.A(databus_out[15]), .B(n33384), .Z(n5_adj_502)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4267_i5_2_lut.init = 16'h2222;
    PFUMX i22680 (.BLUT(n30780), .ALUT(n30779), .C0(\register_addr[1] ), 
          .Z(n30781));
    LUT4 Select_4231_i5_2_lut (.A(databus_out[27]), .B(rw), .Z(n5_adj_574)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4231_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_481 (.A(read_value_adj_309[15]), .B(\read_value[15]_adj_305 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_559)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_481.init = 16'heca0;
    LUT4 i2_4_lut_adj_482 (.A(read_value_adj_309[27]), .B(\read_value[27]_adj_306 ), 
         .C(n52_adj_158), .D(n31446), .Z(n10_adj_575)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_482.init = 16'heca0;
    PWMReceiver recv_ch8 (.GND_net(GND_net), .debug_c_c(debug_c_c), .n33386(n33386), 
            .rc_ch8_c(rc_ch8_c), .n29817(n29817), .n33385(n33385), .\register[6] ({\register[6] }), 
            .n13956(n13956), .n1239(n1239), .n27563(n27563), .n29783(n29783)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(257[14] 261[36])
    PWMReceiver_U1 recv_ch7 (.\register[5] ({\register[5] }), .debug_c_c(debug_c_c), 
            .n33385(n33385), .n33386(n33386), .rc_ch7_c(rc_ch7_c), .GND_net(GND_net), 
            .n33387(n33387), .n1224(n1224), .n27542(n27542), .n29826(n29826)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(252[14] 256[36])
    PWMReceiver_U2 recv_ch4 (.n33385(n33385), .debug_c_c(debug_c_c), .n33386(n33386), 
            .rc_ch4_c(rc_ch4_c), .GND_net(GND_net), .n33387(n33387), .\register[4] ({\register[4] }), 
            .n1209(n1209), .n27549(n27549), .n29837(n29837)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(247[14] 251[36])
    PWMReceiver_U3 recv_ch3 (.debug_c_c(debug_c_c), .n33386(n33386), .rc_ch3_c(rc_ch3_c), 
            .GND_net(GND_net), .n33387(n33387), .\register[3] ({\register[3] }), 
            .n14499(n14499), .n1194(n1194), .n27540(n27540), .n29839(n29839), 
            .n29529(n29529), .n29943(n29943), .n14(n14_adj_307)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(242[14] 246[36])
    PWMReceiver_U4 recv_ch2 (.GND_net(GND_net), .n29831(n29831), .debug_c_c(debug_c_c), 
            .n33386(n33386), .rc_ch2_c(rc_ch2_c), .n31411(n31411), .n33387(n33387), 
            .\register[2] ({\register[2] }), .n14512(n14512), .n29846(n29846), 
            .n1179(n1179), .n27535(n27535), .n33385(n33385), .n31511(n31511)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(237[14] 241[36])
    PWMReceiver_U5 recv_ch1 (.debug_c_c(debug_c_c), .n33386(n33386), .\register[1] ({\register[1] }), 
            .n14513(n14513), .rc_ch1_c(rc_ch1_c), .GND_net(GND_net), .n29829(n29829), 
            .n33385(n33385), .n1164(n1164), .n27546(n27546), .n29810(n29810)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(232[17] 236[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (GND_net, debug_c_c, n33386, rc_ch8_c, n29817, 
            n33385, \register[6] , n13956, n1239, n27563, n29783) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n33386;
    input rc_ch8_c;
    output n29817;
    input n33385;
    output [7:0]\register[6] ;
    input n13956;
    output n1239;
    input n27563;
    output n29783;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n27591, n31466, n31593, n31530, n27755, n31499, n27723, 
        n27394, n10, n26459, n31601;
    wire [15:0]n116;
    
    wire n26460, n31592, n29376, n31479, n1245, n1233, n31542, 
        n26458, n29252, n4, n26457, n26456, n31467, n26455, n29399, 
        n29313, n54, n29553, n23, n28996, n17065, n24;
    wire [7:0]n1137;
    wire [7:0]n43;
    
    wire n31596, n29471, n31531, n29249, n31582, n6, n31594, n4_adj_218, 
        n29400, n26462, n26461, n28987, n29561, n29637, n26734, 
        n26733, n26732, n26731;
    
    LUT4 i15625_2_lut_rep_323 (.A(count[9]), .B(n27591), .Z(n31466)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i15625_2_lut_rep_323.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(count[9]), .B(n27591), .C(n31593), .D(n31530), 
         .Z(n27755)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_4_lut.init = 16'hfff8;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31499), .C(n27723), 
         .D(n27394), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    CCU2D add_1794_11 (.A0(count[9]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31601), .C1(GND_net), .D1(GND_net), .CIN(n26459), 
          .COUT(n26460), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_11.INIT0 = 16'hd222;
    defparam add_1794_11.INIT1 = 16'hd222;
    defparam add_1794_11.INJECT1_0 = "NO";
    defparam add_1794_11.INJECT1_1 = "NO";
    LUT4 i22038_4_lut_rep_336 (.A(n31592), .B(count[13]), .C(count[12]), 
         .D(n29376), .Z(n31479)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i22038_4_lut_rep_336.init = 16'heaaa;
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n33386), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1245));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1245), .SP(n33386), .CK(debug_c_c), .Q(n1233));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_356_4_lut (.A(count[12]), .B(n31592), .C(count[13]), 
         .D(n31542), .Z(n31499)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_356_4_lut.init = 16'hfffe;
    CCU2D add_1794_9 (.A0(count[7]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31601), .C1(GND_net), .D1(GND_net), .CIN(n26458), 
          .COUT(n26459), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_9.INIT0 = 16'hd222;
    defparam add_1794_9.INIT1 = 16'hd222;
    defparam add_1794_9.INJECT1_0 = "NO";
    defparam add_1794_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(count[4]), .B(n31542), .C(n29252), .D(n4), .Z(n29376)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfcec;
    CCU2D add_1794_7 (.A0(count[5]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31601), .C1(GND_net), .D1(GND_net), .CIN(n26457), 
          .COUT(n26458), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_7.INIT0 = 16'hd222;
    defparam add_1794_7.INIT1 = 16'hd222;
    defparam add_1794_7.INJECT1_0 = "NO";
    defparam add_1794_7.INJECT1_1 = "NO";
    CCU2D add_1794_5 (.A0(count[3]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31601), .C1(GND_net), .D1(GND_net), .CIN(n26456), 
          .COUT(n26457), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_5.INIT0 = 16'hd222;
    defparam add_1794_5.INIT1 = 16'hd222;
    defparam add_1794_5.INJECT1_0 = "NO";
    defparam add_1794_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_324_3_lut_4_lut (.A(count[9]), .B(n31593), .C(count[8]), 
         .D(n31530), .Z(n31467)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_324_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_1794_3 (.A0(count[1]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31601), .C1(GND_net), .D1(GND_net), .CIN(n26455), 
          .COUT(n26456), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_3.INIT0 = 16'hd222;
    defparam add_1794_3.INIT1 = 16'hd222;
    defparam add_1794_3.INJECT1_0 = "NO";
    defparam add_1794_3.INJECT1_1 = "NO";
    CCU2D add_1794_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29399), .B1(n1245), .C1(count[0]), .D1(n1233), .COUT(n26455), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_1.INIT0 = 16'hF000;
    defparam add_1794_1.INIT1 = 16'ha565;
    defparam add_1794_1.INJECT1_0 = "NO";
    defparam add_1794_1.INJECT1_1 = "NO";
    LUT4 i21_3_lut_4_lut (.A(n31530), .B(n31542), .C(n27755), .D(n29313), 
         .Z(n54)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i21_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i22357_4_lut (.A(n54), .B(n29553), .C(n23), .D(n10), .Z(n29817)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22357_4_lut.init = 16'h3332;
    LUT4 i3_4_lut (.A(n31592), .B(n28996), .C(n31593), .D(n33385), .Z(n17065)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[13]), .B(n24), .C(count[12]), .D(n29553), 
         .Z(n28996)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i31_3_lut (.A(n29313), .B(n27591), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut (.A(n23), .B(n1137[7]), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_325 (.A(count[8]), .B(n31499), .C(n31596), .D(n29471), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_325.init = 16'h0222;
    LUT4 i1_4_lut_adj_326 (.A(n31596), .B(n31531), .C(count[0]), .D(n29252), 
         .Z(n29313)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_326.init = 16'h8000;
    LUT4 i3_4_lut_adj_327 (.A(count[6]), .B(count[8]), .C(count[7]), .D(n29249), 
         .Z(n27591)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_327.init = 16'hfffe;
    LUT4 i1_4_lut_adj_328 (.A(count[2]), .B(n31582), .C(n6), .D(count[0]), 
         .Z(n29249)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_328.init = 16'hccc8;
    LUT4 i2_2_lut (.A(count[3]), .B(count[1]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i21999_2_lut (.A(n1233), .B(n1245), .Z(n29553)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21999_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_439 (.A(count[4]), .B(count[5]), .Z(n31582)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_439.init = 16'h8888;
    LUT4 i3_4_lut_adj_329 (.A(count[0]), .B(n31594), .C(n31531), .D(n31596), 
         .Z(n27723)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_329.init = 16'h8000;
    LUT4 i2_4_lut (.A(n31594), .B(count[5]), .C(count[4]), .D(n4_adj_218), 
         .Z(n27394)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_2_lut_rep_388_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n31531)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_388_3_lut.init = 16'h8080;
    LUT4 i21919_2_lut_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(n31594), 
         .D(count[3]), .Z(n29471)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i21919_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_330 (.A(n23), .B(n1137[6]), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_330.init = 16'h8888;
    LUT4 i1_2_lut_adj_331 (.A(n23), .B(n1137[5]), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_331.init = 16'h8888;
    LUT4 i1_2_lut_adj_332 (.A(n23), .B(n1137[4]), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_332.init = 16'h8888;
    LUT4 i1_2_lut_adj_333 (.A(n23), .B(n1137[3]), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_333.init = 16'h8888;
    LUT4 i1_2_lut_adj_334 (.A(n23), .B(n1137[2]), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_334.init = 16'h8888;
    LUT4 i22461_3_lut_3_lut_4_lut (.A(n27394), .B(n31467), .C(n27755), 
         .D(n31479), .Z(n29400)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i22461_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_2_lut_adj_335 (.A(n23), .B(n1137[1]), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_335.init = 16'h8888;
    LUT4 i1_2_lut_rep_449 (.A(count[15]), .B(count[14]), .Z(n31592)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_449.init = 16'heeee;
    LUT4 i2_3_lut_rep_387_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n31530)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_387_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_450 (.A(count[11]), .B(count[10]), .Z(n31593)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_450.init = 16'heeee;
    LUT4 i1_2_lut_rep_399_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n31542)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_399_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_451 (.A(count[6]), .B(count[7]), .Z(n31594)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_451.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n29252)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_453 (.A(count[2]), .B(count[1]), .Z(n31596)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_453.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_336 (.A(count[2]), .B(count[1]), .C(count[3]), 
         .Z(n4_adj_218)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_336.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i5_2_lut_rep_458 (.A(n1233), .B(n1245), .Z(n31601)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_458.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_337 (.A(n1233), .B(n1245), .C(n31479), .Z(n29399)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_adj_337.init = 16'hf4f4;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1794_17 (.A0(count[15]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26462), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_17.INIT0 = 16'hd222;
    defparam add_1794_17.INIT1 = 16'h0000;
    defparam add_1794_17.INJECT1_0 = "NO";
    defparam add_1794_17.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13956), .PD(n17065), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX valid_48 (.D(n29400), .SP(n27563), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1239));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_338 (.A(n23), .B(n1137[0]), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_338.init = 16'h8888;
    CCU2D add_1794_15 (.A0(count[13]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31601), .C1(GND_net), .D1(GND_net), .CIN(n26461), 
          .COUT(n26462), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_15.INIT0 = 16'hd222;
    defparam add_1794_15.INIT1 = 16'hd222;
    defparam add_1794_15.INJECT1_0 = "NO";
    defparam add_1794_15.INJECT1_1 = "NO";
    CCU2D add_1794_13 (.A0(count[11]), .B0(n31601), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31601), .C1(GND_net), .D1(GND_net), .CIN(n26460), 
          .COUT(n26461), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1794_13.INIT0 = 16'hd222;
    defparam add_1794_13.INIT1 = 16'hd222;
    defparam add_1794_13.INJECT1_0 = "NO";
    defparam add_1794_13.INJECT1_1 = "NO";
    LUT4 i22323_4_lut (.A(n28987), .B(n31601), .C(n31479), .D(n29553), 
         .Z(n29783)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i22323_4_lut.init = 16'h3031;
    LUT4 i3_4_lut_adj_339 (.A(n31467), .B(n31593), .C(n29561), .D(n29637), 
         .Z(n28987)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_339.init = 16'h0032;
    LUT4 i1_2_lut_adj_340 (.A(n27723), .B(n27394), .Z(n29561)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_340.init = 16'h8888;
    LUT4 i22078_4_lut (.A(n54), .B(n31530), .C(n23), .D(n31466), .Z(n29637)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22078_4_lut.init = 16'hfffe;
    CCU2D sub_78_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26734), 
          .S0(n1137[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_9.INIT1 = 16'h0000;
    defparam sub_78_add_2_9.INJECT1_0 = "NO";
    defparam sub_78_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26733), 
          .COUT(n26734), .S0(n1137[5]), .S1(n1137[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_7.INJECT1_0 = "NO";
    defparam sub_78_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26732), 
          .COUT(n26733), .S0(n1137[3]), .S1(n1137[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_5.INJECT1_0 = "NO";
    defparam sub_78_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26731), 
          .COUT(n26732), .S0(n1137[1]), .S1(n1137[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_3.INJECT1_0 = "NO";
    defparam sub_78_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26731), 
          .S1(n1137[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_1.INIT0 = 16'hF000;
    defparam sub_78_add_2_1.INIT1 = 16'h5555;
    defparam sub_78_add_2_1.INJECT1_0 = "NO";
    defparam sub_78_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (\register[5] , debug_c_c, n33385, n33386, rc_ch7_c, 
            GND_net, n33387, n1224, n27542, n29826) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\register[5] ;
    input debug_c_c;
    input n33385;
    input n33386;
    input rc_ch7_c;
    input GND_net;
    input n33387;
    output n1224;
    input n27542;
    output n29826;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n14450, n16851;
    wire [7:0]n43;
    
    wire n31605, n29607, n54;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n79, n31607, n4, n27302, n1230, n1218, n31603, n31508, 
        n31510, n29280, n13767, n31484, n31606, n31509, n31547, 
        n27714, n31604, n29405, n27588, n31483, n31546, n31452, 
        n29579, n31545, n31451, n29406;
    wire [15:0]n116;
    
    wire n26470, n26469, n26468, n26467, n26466, n13401, n26465, 
        n4_adj_217, n26464, n31485, n26463, n27541, n29629, n26738;
    wire [7:0]n1128;
    
    wire n27614, n6, n26737, n26736, n26735, n28966, n24;
    
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i22335_4_lut_4_lut (.A(n31605), .B(n29607), .C(n33385), .D(n54), 
         .Z(n14450)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22335_4_lut_4_lut.init = 16'h5040;
    LUT4 i1_2_lut (.A(count[5]), .B(count[4]), .Z(n79)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2_4_lut (.A(n31607), .B(count[4]), .C(count[5]), .D(n4), .Z(n27302)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n33386), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1230));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1230), .SP(n33386), .CK(debug_c_c), .Q(n1218));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i21_3_lut_4_lut (.A(n31603), .B(n31508), .C(n31510), .D(n29280), 
         .Z(n54)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i21_3_lut_4_lut.init = 16'h1110;
    LUT4 i1_2_lut_rep_341_3_lut_4_lut (.A(count[9]), .B(n31603), .C(count[8]), 
         .D(n13767), .Z(n31484)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_341_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_366_4_lut (.A(count[3]), .B(n31606), .C(n79), .D(n31607), 
         .Z(n31509)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_366_4_lut.init = 16'h8000;
    LUT4 i5_2_lut_rep_404 (.A(n1218), .B(n1230), .Z(n31547)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_404.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1218), .B(n1230), .C(n27714), .D(n31604), 
         .Z(n29405)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_3_lut_rep_365 (.A(n27588), .B(n13767), .C(count[9]), .Z(n31508)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_3_lut_rep_365.init = 16'hecec;
    LUT4 i2_2_lut_rep_340_4_lut (.A(n27588), .B(n13767), .C(count[9]), 
         .D(n31603), .Z(n31483)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i2_2_lut_rep_340_4_lut.init = 16'hffec;
    LUT4 i1_3_lut_rep_309_4_lut (.A(n31607), .B(n31546), .C(n31510), .D(count[8]), 
         .Z(n31452)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_rep_309_4_lut.init = 16'h0700;
    LUT4 i1_2_lut_3_lut_4_lut_adj_312 (.A(n31607), .B(n31546), .C(n27302), 
         .D(count[0]), .Z(n29579)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut_adj_312.init = 16'h8000;
    LUT4 i1_2_lut_rep_308_3_lut_4_lut (.A(n13767), .B(n31545), .C(n27302), 
         .D(count[8]), .Z(n31451)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_308_3_lut_4_lut.init = 16'hfffe;
    LUT4 i22459_3_lut_3_lut_4_lut (.A(n31604), .B(n27714), .C(n31451), 
         .D(n31483), .Z(n29406)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i22459_3_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    CCU2D add_1790_17 (.A0(count[15]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26470), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_17.INIT0 = 16'hd222;
    defparam add_1790_17.INIT1 = 16'h0000;
    defparam add_1790_17.INJECT1_0 = "NO";
    defparam add_1790_17.INJECT1_1 = "NO";
    CCU2D add_1790_15 (.A0(count[13]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31547), .C1(GND_net), .D1(GND_net), .CIN(n26469), 
          .COUT(n26470), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_15.INIT0 = 16'hd222;
    defparam add_1790_15.INIT1 = 16'hd222;
    defparam add_1790_15.INJECT1_0 = "NO";
    defparam add_1790_15.INJECT1_1 = "NO";
    CCU2D add_1790_13 (.A0(count[11]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31547), .C1(GND_net), .D1(GND_net), .CIN(n26468), 
          .COUT(n26469), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_13.INIT0 = 16'hd222;
    defparam add_1790_13.INIT1 = 16'hd222;
    defparam add_1790_13.INJECT1_0 = "NO";
    defparam add_1790_13.INJECT1_1 = "NO";
    CCU2D add_1790_11 (.A0(count[9]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31547), .C1(GND_net), .D1(GND_net), .CIN(n26467), 
          .COUT(n26468), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_11.INIT0 = 16'hd222;
    defparam add_1790_11.INIT1 = 16'hd222;
    defparam add_1790_11.INJECT1_0 = "NO";
    defparam add_1790_11.INJECT1_1 = "NO";
    CCU2D add_1790_9 (.A0(count[7]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31547), .C1(GND_net), .D1(GND_net), .CIN(n26466), 
          .COUT(n26467), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_9.INIT0 = 16'hd222;
    defparam add_1790_9.INIT1 = 16'hd222;
    defparam add_1790_9.INJECT1_0 = "NO";
    defparam add_1790_9.INJECT1_1 = "NO";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_313 (.A(count[13]), .B(count[12]), .C(n13401), .D(n31545), 
         .Z(n27714)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_313.init = 16'h8880;
    CCU2D add_1790_7 (.A0(count[5]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31547), .C1(GND_net), .D1(GND_net), .CIN(n26465), 
          .COUT(n26466), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_7.INIT0 = 16'hd222;
    defparam add_1790_7.INIT1 = 16'hd222;
    defparam add_1790_7.INJECT1_0 = "NO";
    defparam add_1790_7.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_314 (.A(n31607), .B(count[5]), .C(count[8]), .D(n4_adj_217), 
         .Z(n13401)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_314.init = 16'ha080;
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14450), .PD(n16851), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_460 (.A(count[11]), .B(count[10]), .Z(n31603)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_460.init = 16'heeee;
    LUT4 i1_2_lut_rep_402_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n31545)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_402_3_lut.init = 16'hfefe;
    CCU2D add_1790_5 (.A0(count[3]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31547), .C1(GND_net), .D1(GND_net), .CIN(n26464), 
          .COUT(n26465), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_5.INIT0 = 16'hd222;
    defparam add_1790_5.INIT1 = 16'hd222;
    defparam add_1790_5.INJECT1_0 = "NO";
    defparam add_1790_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_367_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n13767), 
         .D(count[9]), .Z(n31510)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_367_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_461 (.A(count[15]), .B(count[14]), .Z(n31604)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_461.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n13767)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21911_2_lut_rep_462 (.A(n1218), .B(n1230), .Z(n31605)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21911_2_lut_rep_462.init = 16'hdddd;
    LUT4 i3068_2_lut_rep_463 (.A(count[1]), .B(count[2]), .Z(n31606)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3068_2_lut_rep_463.init = 16'h8888;
    LUT4 i3_3_lut_rep_403_4_lut (.A(count[1]), .B(count[2]), .C(n79), 
         .D(count[3]), .Z(n31546)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_3_lut_rep_403_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_217)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_464 (.A(count[7]), .B(count[6]), .Z(n31607)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_464.init = 16'h8888;
    LUT4 i1_2_lut_rep_342_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[0]), 
         .D(n31546), .Z(n31485)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_342_3_lut_4_lut.init = 16'h8000;
    CCU2D add_1790_3 (.A0(count[1]), .B0(n31547), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31547), .C1(GND_net), .D1(GND_net), .CIN(n26463), 
          .COUT(n26464), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_3.INIT0 = 16'hd222;
    defparam add_1790_3.INIT1 = 16'hd222;
    defparam add_1790_3.INJECT1_0 = "NO";
    defparam add_1790_3.INJECT1_1 = "NO";
    CCU2D add_1790_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29405), .B1(n1230), .C1(count[0]), .D1(n1218), .COUT(n26463), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1790_1.INIT0 = 16'hF000;
    defparam add_1790_1.INIT1 = 16'ha565;
    defparam add_1790_1.INJECT1_0 = "NO";
    defparam add_1790_1.INJECT1_1 = "NO";
    FD1P3IX valid_48 (.D(n29406), .SP(n27542), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1224));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i22366_4_lut (.A(n31604), .B(n31547), .C(n27714), .D(n27541), 
         .Z(n29826)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22366_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n31484), .B(n31605), .C(n29629), .D(n29579), .Z(n27541)) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hcfce;
    LUT4 i22070_4_lut (.A(n31603), .B(n54), .C(n31508), .D(n31452), 
         .Z(n29629)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22070_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_315 (.A(n31546), .B(n31607), .C(count[8]), .D(count[0]), 
         .Z(n29280)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_315.init = 16'h8000;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    CCU2D sub_77_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26738), 
          .S0(n1128[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_9.INIT1 = 16'h0000;
    defparam sub_77_add_2_9.INJECT1_0 = "NO";
    defparam sub_77_add_2_9.INJECT1_1 = "NO";
    LUT4 i3_4_lut (.A(n27614), .B(n6), .C(count[8]), .D(n79), .Z(n27588)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_4_lut.init = 16'hfefc;
    CCU2D sub_77_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26737), 
          .COUT(n26738), .S0(n1128[5]), .S1(n1128[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_7.INJECT1_0 = "NO";
    defparam sub_77_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26736), 
          .COUT(n26737), .S0(n1128[3]), .S1(n1128[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_5.INJECT1_0 = "NO";
    defparam sub_77_add_2_5.INJECT1_1 = "NO";
    LUT4 i22048_4_lut_4_lut (.A(n27302), .B(n31484), .C(n31485), .D(n31452), 
         .Z(n29607)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;
    defparam i22048_4_lut_4_lut.init = 16'hff02;
    LUT4 i1_2_lut_4_lut (.A(count[8]), .B(n31509), .C(n31510), .D(n1128[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0200;
    CCU2D sub_77_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26735), 
          .COUT(n26736), .S0(n1128[1]), .S1(n1128[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_3.INJECT1_0 = "NO";
    defparam sub_77_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_316 (.A(count[8]), .B(n31509), .C(n31510), 
         .D(n1128[1]), .Z(n43[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_316.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_317 (.A(count[8]), .B(n31509), .C(n31510), 
         .D(n1128[4]), .Z(n43[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_317.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_318 (.A(count[8]), .B(n31509), .C(n31510), 
         .D(n1128[5]), .Z(n43[5])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_318.init = 16'h0200;
    CCU2D sub_77_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26735), 
          .S1(n1128[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_1.INIT0 = 16'hF000;
    defparam sub_77_add_2_1.INIT1 = 16'h5555;
    defparam sub_77_add_2_1.INJECT1_0 = "NO";
    defparam sub_77_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_319 (.A(count[8]), .B(n31509), .C(n31510), 
         .D(n1128[6]), .Z(n43[6])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_319.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_320 (.A(count[8]), .B(n31509), .C(n31510), 
         .D(n1128[7]), .Z(n43[7])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_320.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_321 (.A(count[8]), .B(n31509), .C(n31510), 
         .D(n1128[0]), .Z(n43[0])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_321.init = 16'h0200;
    LUT4 i3_4_lut_adj_322 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27614)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_322.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_323 (.A(count[8]), .B(n31509), .C(n31510), 
         .D(n1128[2]), .Z(n43[2])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_323.init = 16'h0200;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_324 (.A(n31604), .B(n28966), .C(n31603), .D(n33385), 
         .Z(n16851)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_324.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[13]), .B(n24), .C(count[12]), .D(n31605), 
         .Z(n28966)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i31_3_lut (.A(n29280), .B(n27588), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (n33385, debug_c_c, n33386, rc_ch4_c, GND_net, 
            n33387, \register[4] , n1209, n27549, n29837) /* synthesis syn_module_defined=1 */ ;
    input n33385;
    input debug_c_c;
    input n33386;
    input rc_ch4_c;
    input GND_net;
    input n33387;
    output [7:0]\register[4] ;
    output n1209;
    input n27549;
    output n29837;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31558, n31516, n29290, n31557, n124, n31488, n31554, 
        n4, n31432, n14490, n31556, n27644, n31433, n22310, n29315, 
        n1215, n1203, n31489, n31455, n5, n27365, n31454, n29304, 
        n13676, n5_adj_212, n29316, n4_adj_213, n4_adj_214, n31515, 
        n31559, n29643, n31563, n103, n26478;
    wire [15:0]n116;
    
    wire n26477, n26476, n26475, n152, n154, n16890;
    wire [7:0]n43;
    
    wire n26474, n26473, n26472, n26471, n6, n29576, n4_adj_216;
    wire [7:0]n1119;
    
    wire n11, n8, n27547, n26742, n26741, n26740, n26739;
    
    LUT4 i1_3_lut_4_lut (.A(count[8]), .B(n31558), .C(count[0]), .D(n31516), 
         .Z(n29290)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_345_4_lut (.A(count[3]), .B(n31557), .C(n124), .D(n31558), 
         .Z(n31488)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_345_4_lut.init = 16'h8000;
    LUT4 i22487_4_lut_4_lut (.A(n31554), .B(n4), .C(n33385), .D(n31432), 
         .Z(n14490)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22487_4_lut_4_lut.init = 16'h5010;
    LUT4 i22454_3_lut_3_lut_4_lut (.A(n31556), .B(n27644), .C(n31433), 
         .D(n22310), .Z(n29315)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i22454_3_lut_3_lut_4_lut.init = 16'h0010;
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n33386), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1215));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1215), .SP(n33386), .CK(debug_c_c), .Q(n1203));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n29290), .B(n22310), .C(n31489), .D(n31455), 
         .Z(n5)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    LUT4 i1_4_lut_4_lut (.A(n27365), .B(n31454), .C(n29304), .D(n31455), 
         .Z(n4)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i1_4_lut_4_lut.init = 16'hfd00;
    LUT4 i1_3_lut_rep_312_4_lut (.A(n31558), .B(n31516), .C(count[8]), 
         .D(n31489), .Z(n31455)) /* synthesis lut_function=(A (B+((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1_3_lut_rep_312_4_lut.init = 16'hff8f;
    LUT4 i1_2_lut_rep_346 (.A(count[9]), .B(n13676), .Z(n31489)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_346.init = 16'heeee;
    LUT4 i1_2_lut_rep_311_3_lut (.A(count[9]), .B(n13676), .C(count[8]), 
         .Z(n31454)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_311_3_lut.init = 16'hfefe;
    LUT4 i21_3_lut_rep_289_4_lut (.A(count[9]), .B(n13676), .C(n22310), 
         .D(n29290), .Z(n31432)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i21_3_lut_rep_289_4_lut.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_290_3_lut_4_lut (.A(count[9]), .B(n13676), .C(n27365), 
         .D(count[8]), .Z(n31433)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_290_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_411 (.A(n1215), .B(n1203), .Z(n31554)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_411.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_413 (.A(count[15]), .B(count[14]), .Z(n31556)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_413.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5_adj_212), 
         .D(n27644), .Z(n29316)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_414 (.A(count[2]), .B(count[1]), .Z(n31557)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_414.init = 16'h8888;
    LUT4 i1_3_lut_rep_373_4_lut (.A(count[2]), .B(count[1]), .C(n124), 
         .D(count[3]), .Z(n31516)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_rep_373_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4_adj_213)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut_adj_305 (.A(count[2]), .B(count[1]), .C(count[5]), 
         .D(count[3]), .Z(n4_adj_214)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut_adj_305.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_415 (.A(count[7]), .B(count[6]), .Z(n31558)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_415.init = 16'h8888;
    LUT4 i1_2_lut_rep_372_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n31515)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_372_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_306 (.A(count[7]), .B(count[6]), .C(count[0]), 
         .D(n31516), .Z(n29304)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut_adj_306.init = 16'h8000;
    LUT4 i21935_2_lut_rep_416 (.A(count[11]), .B(count[10]), .Z(n31559)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21935_2_lut_rep_416.init = 16'heeee;
    LUT4 i22084_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n29643)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22084_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_420 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n31563)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_420.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_307 (.A(count[7]), .B(count[6]), .C(count[8]), 
         .D(n124), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_307.init = 16'hfffe;
    CCU2D add_1786_17 (.A0(count[15]), .B0(n5_adj_212), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26478), .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_17.INIT0 = 16'hd222;
    defparam add_1786_17.INIT1 = 16'h0000;
    defparam add_1786_17.INJECT1_0 = "NO";
    defparam add_1786_17.INJECT1_1 = "NO";
    CCU2D add_1786_15 (.A0(count[13]), .B0(n5_adj_212), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n5_adj_212), .C1(GND_net), 
          .D1(GND_net), .CIN(n26477), .COUT(n26478), .S0(n116[13]), 
          .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_15.INIT0 = 16'hd222;
    defparam add_1786_15.INIT1 = 16'hd222;
    defparam add_1786_15.INJECT1_0 = "NO";
    defparam add_1786_15.INJECT1_1 = "NO";
    CCU2D add_1786_13 (.A0(count[11]), .B0(n5_adj_212), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n5_adj_212), .C1(GND_net), 
          .D1(GND_net), .CIN(n26476), .COUT(n26477), .S0(n116[11]), 
          .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_13.INIT0 = 16'hd222;
    defparam add_1786_13.INIT1 = 16'hd222;
    defparam add_1786_13.INJECT1_0 = "NO";
    defparam add_1786_13.INJECT1_1 = "NO";
    CCU2D add_1786_11 (.A0(count[9]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26475), .COUT(n26476), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_11.INIT0 = 16'hd222;
    defparam add_1786_11.INIT1 = 16'hd222;
    defparam add_1786_11.INJECT1_0 = "NO";
    defparam add_1786_11.INJECT1_1 = "NO";
    PFUMX i14065 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    CCU2D add_1786_9 (.A0(count[7]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26474), .COUT(n26475), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_9.INIT0 = 16'hd222;
    defparam add_1786_9.INIT1 = 16'hd222;
    defparam add_1786_9.INJECT1_0 = "NO";
    defparam add_1786_9.INJECT1_1 = "NO";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1786_7 (.A0(count[5]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26473), .COUT(n26474), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_7.INIT0 = 16'hd222;
    defparam add_1786_7.INIT1 = 16'hd222;
    defparam add_1786_7.INJECT1_0 = "NO";
    defparam add_1786_7.INJECT1_1 = "NO";
    CCU2D add_1786_5 (.A0(count[3]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26472), .COUT(n26473), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_5.INIT0 = 16'hd222;
    defparam add_1786_5.INIT1 = 16'hd222;
    defparam add_1786_5.INJECT1_0 = "NO";
    defparam add_1786_5.INJECT1_1 = "NO";
    CCU2D add_1786_3 (.A0(count[1]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26471), .COUT(n26472), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_3.INIT0 = 16'hd222;
    defparam add_1786_3.INIT1 = 16'hd222;
    defparam add_1786_3.INJECT1_0 = "NO";
    defparam add_1786_3.INJECT1_1 = "NO";
    CCU2D add_1786_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29316), .B1(n1215), .C1(count[0]), .D1(n1203), .COUT(n26471), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1786_1.INIT0 = 16'hF000;
    defparam add_1786_1.INIT1 = 16'ha565;
    defparam add_1786_1.INJECT1_0 = "NO";
    defparam add_1786_1.INJECT1_1 = "NO";
    LUT4 i23_4_lut (.A(n31563), .B(count[2]), .C(n124), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(count[4]), .B(count[5]), .Z(n124)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i22019_3_lut_4_lut (.A(count[8]), .B(n31489), .C(n27365), .D(n29304), 
         .Z(n29576)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22019_3_lut_4_lut.init = 16'hfeee;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n31559), .D(n4_adj_216), 
         .Z(n27644)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut (.A(count[9]), .B(count[4]), .C(n31515), .D(n4_adj_214), 
         .Z(n4_adj_216)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfaea;
    LUT4 i15416_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15416_2_lut_4_lut.init = 16'h0400;
    LUT4 i2_4_lut_adj_308 (.A(n33385), .B(n31556), .C(n11), .D(n29643), 
         .Z(n16890)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_308.init = 16'h0020;
    LUT4 i15415_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15415_2_lut_4_lut.init = 16'h0400;
    LUT4 i15414_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15414_2_lut_4_lut.init = 16'h0400;
    LUT4 i4_4_lut (.A(n29290), .B(n8), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0c88;
    FD1P3IX valid_48 (.D(n29315), .SP(n27549), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1209));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i22377_4_lut (.A(n31556), .B(n5_adj_212), .C(n27644), .D(n27547), 
         .Z(n29837)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22377_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_309 (.A(n5), .B(n31554), .C(n29576), .D(n22310), 
         .Z(n27547)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_309.init = 16'hccec;
    LUT4 i15413_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15413_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_adj_310 (.A(n1203), .B(n1215), .Z(n8)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_adj_310.init = 16'h2222;
    LUT4 i15412_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15412_2_lut_4_lut.init = 16'h0400;
    LUT4 i15411_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15411_2_lut_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14490), .PD(n16890), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i15410_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15410_2_lut_4_lut.init = 16'h0400;
    LUT4 i15196_2_lut_4_lut (.A(n31489), .B(count[8]), .C(n31488), .D(n1119[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15196_2_lut_4_lut.init = 16'h0400;
    CCU2D sub_76_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26742), 
          .S0(n1119[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_9.INIT1 = 16'h0000;
    defparam sub_76_add_2_9.INJECT1_0 = "NO";
    defparam sub_76_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26741), 
          .COUT(n26742), .S0(n1119[5]), .S1(n1119[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_7.INJECT1_0 = "NO";
    defparam sub_76_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26740), 
          .COUT(n26741), .S0(n1119[3]), .S1(n1119[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_5.INJECT1_0 = "NO";
    defparam sub_76_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26739), 
          .COUT(n26740), .S0(n1119[1]), .S1(n1119[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_3.INJECT1_0 = "NO";
    defparam sub_76_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26739), 
          .S1(n1119[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_1.INIT0 = 16'hF000;
    defparam sub_76_add_2_1.INIT1 = 16'h5555;
    defparam sub_76_add_2_1.INJECT1_0 = "NO";
    defparam sub_76_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_311 (.A(n31558), .B(count[5]), .C(count[3]), .D(n4_adj_213), 
         .Z(n27365)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_311.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n31556), .D(n31559), 
         .Z(n13676)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(n1203), .B(n1215), .Z(n5_adj_212)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i15574_3_lut (.A(count[9]), .B(n13676), .C(n154), .Z(n22310)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15574_3_lut.init = 16'hecec;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (debug_c_c, n33386, rc_ch3_c, GND_net, n33387, 
            \register[3] , n14499, n1194, n27540, n29839, n29529, 
            n29943, n14) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n33386;
    input rc_ch3_c;
    input GND_net;
    input n33387;
    output [7:0]\register[3] ;
    input n14499;
    output n1194;
    input n27540;
    output n29839;
    output n29529;
    output n29943;
    input n14;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n1188, n1200, n5;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31564, n31571, n31573, n31492, n26486;
    wire [15:0]n116;
    
    wire n26485, n13662, n31491, n31457, n31458, n31521, n29301, 
        n27277, n29591, n31438, n29409, n26484, n154, n26483, 
        n31561, n103, n26482, n5_adj_208, n54, n7, n6, n31524, 
        n4, n4_adj_209, n31574, n27716, n29408, n26481, n26480, 
        n26479;
    wire [7:0]n1110;
    wire [7:0]n43;
    
    wire n16900, n152, n6_adj_210, n27539, n29594, n26746, n26745, 
        n26744, n26743, n29343, n4_adj_211, n10, n29649, n26;
    
    LUT4 i5_2_lut (.A(n1188), .B(n1200), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i3_3_lut_rep_349_4_lut (.A(count[3]), .B(n31564), .C(n31571), 
         .D(n31573), .Z(n31492)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_3_lut_rep_349_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n33386), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1200));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1200), .SP(n33386), .CK(debug_c_c), .Q(n1188));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D add_1782_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26486), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_17.INIT0 = 16'hd222;
    defparam add_1782_17.INIT1 = 16'h0000;
    defparam add_1782_17.INJECT1_0 = "NO";
    defparam add_1782_17.INJECT1_1 = "NO";
    CCU2D add_1782_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26485), 
          .COUT(n26486), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_15.INIT0 = 16'hd222;
    defparam add_1782_15.INIT1 = 16'hd222;
    defparam add_1782_15.INJECT1_0 = "NO";
    defparam add_1782_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_348 (.A(count[9]), .B(n13662), .Z(n31491)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_348.init = 16'heeee;
    LUT4 i1_2_lut_rep_314_3_lut (.A(count[9]), .B(n13662), .C(count[8]), 
         .Z(n31457)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_314_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_315_4_lut (.A(count[9]), .B(n13662), .C(n31492), 
         .D(count[8]), .Z(n31458)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i2_3_lut_rep_315_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_4_lut (.A(n31573), .B(n31571), .C(n31521), .D(count[0]), 
         .Z(n29301)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i22452_3_lut_3_lut_4_lut (.A(n27277), .B(n31457), .C(n29591), 
         .D(n31438), .Z(n29409)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i22452_3_lut_3_lut_4_lut.init = 16'h000e;
    CCU2D add_1782_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26484), 
          .COUT(n26485), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_13.INIT0 = 16'hd222;
    defparam add_1782_13.INIT1 = 16'hd222;
    defparam add_1782_13.INJECT1_0 = "NO";
    defparam add_1782_13.INJECT1_1 = "NO";
    LUT4 i22033_3_lut (.A(n13662), .B(count[9]), .C(n154), .Z(n29591)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i22033_3_lut.init = 16'heaea;
    CCU2D add_1782_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26483), 
          .COUT(n26484), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_11.INIT0 = 16'hd222;
    defparam add_1782_11.INIT1 = 16'hd222;
    defparam add_1782_11.INJECT1_0 = "NO";
    defparam add_1782_11.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_418 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n31561)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_418.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_300 (.A(count[7]), .B(count[6]), .C(count[8]), 
         .D(n31564), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_300.init = 16'hfffe;
    CCU2D add_1782_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26482), 
          .COUT(n26483), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_9.INIT0 = 16'hd222;
    defparam add_1782_9.INIT1 = 16'hd222;
    defparam add_1782_9.INJECT1_0 = "NO";
    defparam add_1782_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_421 (.A(count[4]), .B(count[5]), .Z(n31564)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_421.init = 16'h8888;
    LUT4 i1_2_lut_rep_378_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n31521)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_378_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n5_adj_208)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_428 (.A(count[7]), .B(count[6]), .Z(n31571)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_428.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_301 (.A(n31491), .B(count[8]), .C(n31492), 
         .D(n54), .Z(n7)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_301.init = 16'h00fb;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n31573), 
         .D(count[8]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_381_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n31524)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_381_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_430 (.A(count[2]), .B(count[1]), .Z(n31573)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_430.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4_adj_209)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_431 (.A(count[15]), .B(count[14]), .Z(n31574)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_431.init = 16'heeee;
    LUT4 i1_2_lut_rep_295_3_lut (.A(count[15]), .B(count[14]), .C(n27716), 
         .Z(n31438)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_295_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_302 (.A(count[15]), .B(count[14]), .C(n5), 
         .D(n27716), .Z(n29408)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_302.init = 16'hfffe;
    CCU2D add_1782_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26481), 
          .COUT(n26482), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_7.INIT0 = 16'hd222;
    defparam add_1782_7.INIT1 = 16'hd222;
    defparam add_1782_7.INJECT1_0 = "NO";
    defparam add_1782_7.INJECT1_1 = "NO";
    CCU2D add_1782_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26480), 
          .COUT(n26481), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_5.INIT0 = 16'hd222;
    defparam add_1782_5.INIT1 = 16'hd222;
    defparam add_1782_5.INJECT1_0 = "NO";
    defparam add_1782_5.INJECT1_1 = "NO";
    CCU2D add_1782_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26479), 
          .COUT(n26480), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_3.INIT0 = 16'hd222;
    defparam add_1782_3.INIT1 = 16'hd222;
    defparam add_1782_3.INJECT1_0 = "NO";
    defparam add_1782_3.INJECT1_1 = "NO";
    CCU2D add_1782_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29408), .B1(n1200), .C1(count[0]), .D1(n1188), .COUT(n26479), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1782_1.INIT0 = 16'hF000;
    defparam add_1782_1.INIT1 = 16'ha565;
    defparam add_1782_1.INJECT1_0 = "NO";
    defparam add_1782_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    LUT4 i15184_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15184_2_lut_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    PFUMX i14314 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i23_4_lut (.A(n31561), .B(count[2]), .C(n31564), .D(n6_adj_210), 
         .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6_adj_210)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3IX valid_48 (.D(n29409), .SP(n27540), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1194));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i22379_4_lut (.A(n31574), .B(n5), .C(n27716), .D(n27539), .Z(n29839)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22379_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n29591), .B(n29529), .C(n7), .D(n29594), .Z(n27539)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14499), .PD(n16900), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D sub_75_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26746), 
          .S0(n1110[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_9.INIT1 = 16'h0000;
    defparam sub_75_add_2_9.INJECT1_0 = "NO";
    defparam sub_75_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26745), 
          .COUT(n26746), .S0(n1110[5]), .S1(n1110[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_7.INJECT1_0 = "NO";
    defparam sub_75_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26744), 
          .COUT(n26745), .S0(n1110[3]), .S1(n1110[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_5.INJECT1_0 = "NO";
    defparam sub_75_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26743), 
          .COUT(n26744), .S0(n1110[1]), .S1(n1110[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_3.INJECT1_0 = "NO";
    defparam sub_75_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26743), 
          .S1(n1110[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_1.INIT0 = 16'hF000;
    defparam sub_75_add_2_1.INIT1 = 16'h5555;
    defparam sub_75_add_2_1.INJECT1_0 = "NO";
    defparam sub_75_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n29343), .D(n4_adj_211), 
         .Z(n27716)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_303 (.A(count[9]), .B(count[4]), .C(n31524), .D(n4_adj_209), 
         .Z(n4_adj_211)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_303.init = 16'hfaea;
    LUT4 i1_2_lut (.A(count[10]), .B(count[11]), .Z(n29343)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31491), .C(n29301), 
         .D(n27277), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22035_3_lut_4_lut (.A(count[8]), .B(n31491), .C(n27277), .D(n29301), 
         .Z(n29594)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22035_3_lut_4_lut.init = 16'hfeee;
    LUT4 i15409_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15409_2_lut_4_lut.init = 16'h0400;
    LUT4 i15408_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15408_2_lut_4_lut.init = 16'h0400;
    LUT4 i15407_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15407_2_lut_4_lut.init = 16'h0400;
    LUT4 i15406_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15406_2_lut_4_lut.init = 16'h0400;
    LUT4 i22483_4_lut (.A(n54), .B(n29529), .C(n31458), .D(n10), .Z(n29943)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22483_4_lut.init = 16'h3323;
    LUT4 i15405_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15405_2_lut_4_lut.init = 16'h0400;
    LUT4 i8_4_lut (.A(n29649), .B(count[10]), .C(n14), .D(n26), .Z(n16900)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i8_4_lut.init = 16'h1000;
    LUT4 i22090_4_lut (.A(count[12]), .B(count[13]), .C(count[11]), .D(n31574), 
         .Z(n29649)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22090_4_lut.init = 16'hfffe;
    LUT4 i33_4_lut (.A(count[8]), .B(n154), .C(count[9]), .D(n29301), 
         .Z(n26)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_4_lut.init = 16'h3a30;
    LUT4 i15404_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15404_2_lut_4_lut.init = 16'h0400;
    LUT4 i15403_2_lut_4_lut (.A(n31491), .B(count[8]), .C(n31492), .D(n1110[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15403_2_lut_4_lut.init = 16'h0400;
    LUT4 i21975_2_lut (.A(n1188), .B(n1200), .Z(n29529)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21975_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_adj_304 (.A(n31571), .B(count[5]), .C(count[3]), .D(n4), 
         .Z(n27277)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_304.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(n31574), .C(count[13]), .D(n29343), 
         .Z(n13662)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(n5_adj_208), .B(n29591), .C(n31491), .D(n6), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (GND_net, n29831, debug_c_c, n33386, rc_ch2_c, 
            n31411, n33387, \register[2] , n14512, n29846, n1179, 
            n27535, n33385, n31511) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n29831;
    input debug_c_c;
    input n33386;
    input rc_ch2_c;
    input n31411;
    input n33387;
    output [7:0]\register[2] ;
    input n14512;
    output n29846;
    output n1179;
    input n27535;
    input n33385;
    input n31511;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26490;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31572;
    wire [15:0]n116;
    
    wire n26491, n29350, n27564, n4, n29351, n29186, n26489, n13701, 
        n26488, n26487, n31481, n29396, n1185, n1173, n13630, 
        n31493, n31459, n31494, n22409, n27661, n31436, n129_adj_206, 
        n31460, n29517, n23, n29653, n29397, n31565, n27608, n31569, 
        n31598, n16909;
    wire [7:0]n43;
    
    wire n31437, n18, n29247, n26494, n26750;
    wire [7:0]n1101;
    
    wire n26749, n26748, n26747, n28998, n4_adj_207, n5, n6, n27517, 
        n26493, n26492;
    
    CCU2D add_1778_9 (.A0(count[7]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31572), .C1(GND_net), .D1(GND_net), .CIN(n26490), 
          .COUT(n26491), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_9.INIT0 = 16'hd222;
    defparam add_1778_9.INIT1 = 16'hd222;
    defparam add_1778_9.INJECT1_0 = "NO";
    defparam add_1778_9.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n29350), .B(count[9]), .C(n27564), .D(n4), .Z(n29351)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut.init = 16'hfeee;
    LUT4 i2_4_lut_adj_288 (.A(count[1]), .B(count[5]), .C(n29186), .D(count[4]), 
         .Z(n27564)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_288.init = 16'hffec;
    LUT4 i1_2_lut (.A(count[10]), .B(count[11]), .Z(n29350)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_289 (.A(count[3]), .B(count[2]), .Z(n29186)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_289.init = 16'h8888;
    CCU2D add_1778_7 (.A0(count[5]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31572), .C1(GND_net), .D1(GND_net), .CIN(n26489), 
          .COUT(n26490), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_7.INIT0 = 16'hd222;
    defparam add_1778_7.INIT1 = 16'hd222;
    defparam add_1778_7.INJECT1_0 = "NO";
    defparam add_1778_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_290 (.A(count[15]), .B(count[14]), .Z(n13701)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_290.init = 16'heeee;
    CCU2D add_1778_5 (.A0(count[3]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31572), .C1(GND_net), .D1(GND_net), .CIN(n26488), 
          .COUT(n26489), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_5.INIT0 = 16'hd222;
    defparam add_1778_5.INIT1 = 16'hd222;
    defparam add_1778_5.INJECT1_0 = "NO";
    defparam add_1778_5.INJECT1_1 = "NO";
    CCU2D add_1778_3 (.A0(count[1]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31572), .C1(GND_net), .D1(GND_net), .CIN(n26487), 
          .COUT(n26488), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_3.INIT0 = 16'hd222;
    defparam add_1778_3.INIT1 = 16'hd222;
    defparam add_1778_3.INJECT1_0 = "NO";
    defparam add_1778_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_338 (.A(n13701), .B(count[13]), .C(count[12]), .D(n29351), 
         .Z(n31481)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_338.init = 16'heaaa;
    CCU2D add_1778_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29396), .B1(n1185), .C1(count[0]), .D1(n1173), .COUT(n26487), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_1.INIT0 = 16'hF000;
    defparam add_1778_1.INIT1 = 16'ha565;
    defparam add_1778_1.INJECT1_0 = "NO";
    defparam add_1778_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_350 (.A(count[9]), .B(n13630), .Z(n31493)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_350.init = 16'heeee;
    LUT4 i1_2_lut_rep_316_3_lut (.A(count[9]), .B(n13630), .C(count[8]), 
         .Z(n31459)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_316_3_lut.init = 16'hfefe;
    LUT4 i15666_2_lut_3_lut_4_lut (.A(count[9]), .B(n13630), .C(n31494), 
         .D(count[8]), .Z(n22409)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i15666_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_293_3_lut_4_lut (.A(count[9]), .B(n13630), .C(n27661), 
         .D(count[8]), .Z(n31436)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_293_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_351 (.A(n129_adj_206), .B(count[1]), .C(count[0]), 
         .Z(n31494)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_3_lut_rep_351.init = 16'h8080;
    LUT4 i1_2_lut_rep_317_4_lut (.A(n129_adj_206), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n31460)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_317_4_lut.init = 16'h8000;
    LUT4 i22094_3_lut_4_lut (.A(n31460), .B(n29517), .C(n31493), .D(n23), 
         .Z(n29653)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i22094_3_lut_4_lut.init = 16'hfffe;
    LUT4 i22447_3_lut_4_lut_4_lut (.A(n31481), .B(n29517), .C(n31459), 
         .D(n27661), .Z(n29397)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i22447_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i1_2_lut_rep_422 (.A(n1185), .B(n1173), .Z(n31565)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_422.init = 16'hbbbb;
    LUT4 i22371_2_lut_3_lut (.A(n1185), .B(n1173), .C(n27608), .Z(n29831)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i22371_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_426 (.A(count[5]), .B(count[4]), .Z(n31569)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_426.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(count[5]), .B(count[4]), .C(n29186), .D(n31598), 
         .Z(n129_adj_206)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n33386), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1185));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i5_2_lut_rep_429 (.A(n1173), .B(n1185), .Z(n31572)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_429.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n1173), .B(n1185), .C(n31481), .Z(n29396)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31411), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31411), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31411), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31411), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31411), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31411), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31411), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31411), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1185), .SP(n33386), .CK(debug_c_c), .Q(n1173));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i21_3_lut_rep_294_4_lut (.A(count[8]), .B(n31494), .C(n31493), 
         .D(n29517), .Z(n31437)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21_3_lut_rep_294_4_lut.init = 16'h00f8;
    LUT4 i1_2_lut_3_lut_adj_291 (.A(count[8]), .B(n31494), .C(count[9]), 
         .Z(n18)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_291.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_455 (.A(count[6]), .B(count[7]), .Z(n31598)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_455.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_292 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_adj_292.init = 16'h8080;
    LUT4 i22386_4_lut (.A(n29247), .B(n31572), .C(n31481), .D(n31565), 
         .Z(n29846)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i22386_4_lut.init = 16'h3031;
    LUT4 i3_4_lut (.A(n31459), .B(n29653), .C(n31494), .D(n27661), .Z(n29247)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut.init = 16'h3222;
    FD1P3IX valid_48 (.D(n29397), .SP(n27535), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1179));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D add_1778_17 (.A0(count[15]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26494), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_17.INIT0 = 16'hd222;
    defparam add_1778_17.INIT1 = 16'h0000;
    defparam add_1778_17.INJECT1_0 = "NO";
    defparam add_1778_17.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26750), 
          .S0(n1101[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_9.INIT1 = 16'h0000;
    defparam sub_74_add_2_9.INJECT1_0 = "NO";
    defparam sub_74_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26749), 
          .COUT(n26750), .S0(n1101[5]), .S1(n1101[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_7.INJECT1_0 = "NO";
    defparam sub_74_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26748), 
          .COUT(n26749), .S0(n1101[3]), .S1(n1101[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_5.INJECT1_0 = "NO";
    defparam sub_74_add_2_5.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14512), .PD(n16909), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D sub_74_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26747), 
          .COUT(n26748), .S0(n1101[1]), .S1(n1101[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_3.INJECT1_0 = "NO";
    defparam sub_74_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26747), 
          .S1(n1101[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_1.INIT0 = 16'hF000;
    defparam sub_74_add_2_1.INIT1 = 16'h5555;
    defparam sub_74_add_2_1.INJECT1_0 = "NO";
    defparam sub_74_add_2_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_293 (.A(n33385), .B(n28998), .C(n1173), .D(n29517), 
         .Z(n16909)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_293.init = 16'h0080;
    LUT4 i3_4_lut_adj_294 (.A(n27608), .B(n1185), .C(n31511), .D(n18), 
         .Z(n28998)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_294.init = 16'h0200;
    LUT4 i15402_2_lut (.A(n1101[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15402_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(count[8]), .B(n31493), .C(count[1]), .D(n129_adj_206), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0222;
    LUT4 i2_4_lut_adj_295 (.A(n31437), .B(n23), .C(n31436), .D(n22409), 
         .Z(n27608)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_295.init = 16'heefe;
    LUT4 i2_4_lut_adj_296 (.A(n31598), .B(count[4]), .C(count[5]), .D(n4_adj_207), 
         .Z(n27661)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_296.init = 16'ha080;
    LUT4 i1_3_lut (.A(count[3]), .B(count[1]), .C(count[2]), .Z(n4_adj_207)) /* synthesis lut_function=(A+(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut.init = 16'heaea;
    LUT4 i21963_4_lut (.A(n13630), .B(count[9]), .C(n5), .D(n6), .Z(n29517)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i21963_4_lut.init = 16'heeea;
    LUT4 i1_2_lut_adj_297 (.A(count[8]), .B(count[6]), .Z(n5)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_adj_297.init = 16'heeee;
    LUT4 i2_4_lut_adj_298 (.A(count[7]), .B(count[3]), .C(n31569), .D(n27517), 
         .Z(n6)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i2_4_lut_adj_298.init = 16'hfaea;
    LUT4 i2_3_lut (.A(count[0]), .B(count[2]), .C(count[1]), .Z(n27517)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i3_4_lut_adj_299 (.A(count[12]), .B(count[13]), .C(n13701), .D(n29350), 
         .Z(n13630)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_299.init = 16'hfffe;
    LUT4 i15401_2_lut (.A(n1101[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15401_2_lut.init = 16'h8888;
    LUT4 i15400_2_lut (.A(n1101[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15400_2_lut.init = 16'h8888;
    LUT4 i15399_2_lut (.A(n1101[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15399_2_lut.init = 16'h8888;
    LUT4 i15398_2_lut (.A(n1101[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15398_2_lut.init = 16'h8888;
    LUT4 i15397_2_lut (.A(n1101[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15397_2_lut.init = 16'h8888;
    LUT4 i15396_2_lut (.A(n1101[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15396_2_lut.init = 16'h8888;
    LUT4 i15175_2_lut (.A(n1101[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15175_2_lut.init = 16'h8888;
    CCU2D add_1778_15 (.A0(count[13]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31572), .C1(GND_net), .D1(GND_net), .CIN(n26493), 
          .COUT(n26494), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_15.INIT0 = 16'hd222;
    defparam add_1778_15.INIT1 = 16'hd222;
    defparam add_1778_15.INJECT1_0 = "NO";
    defparam add_1778_15.INJECT1_1 = "NO";
    CCU2D add_1778_13 (.A0(count[11]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31572), .C1(GND_net), .D1(GND_net), .CIN(n26492), 
          .COUT(n26493), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_13.INIT0 = 16'hd222;
    defparam add_1778_13.INIT1 = 16'hd222;
    defparam add_1778_13.INJECT1_0 = "NO";
    defparam add_1778_13.INJECT1_1 = "NO";
    CCU2D add_1778_11 (.A0(count[9]), .B0(n31572), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31572), .C1(GND_net), .D1(GND_net), .CIN(n26491), 
          .COUT(n26492), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_11.INIT0 = 16'hd222;
    defparam add_1778_11.INIT1 = 16'hd222;
    defparam add_1778_11.INJECT1_0 = "NO";
    defparam add_1778_11.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (debug_c_c, n33386, \register[1] , n14513, rc_ch1_c, 
            GND_net, n29829, n33385, n1164, n27546, n29810) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n33386;
    output [7:0]\register[1] ;
    input n14513;
    input rc_ch1_c;
    input GND_net;
    output n29829;
    input n33385;
    output n1164;
    input n27546;
    output n29810;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31576, n29365, n31495, n31578, n31579, n31577, n29286, 
        n1158, n1170, n29110, n31441, n33381, n31439, n29402, 
        n27607, n10, n31440, n31527, n31461, n28947, n7, n10_adj_204, 
        n29568, n27647, n16912;
    wire [7:0]n43;
    
    wire n5, n29403, n31528, n29109, n31526, n26502;
    wire [15:0]n116;
    
    wire n26501, n26500, n29523, n26499, n26498, n16, n26, n26497;
    wire [7:0]n1092;
    
    wire n26754, n26753, n27574, n6, n26496, n26495, n26752, n26751, 
        n6_adj_205, n4, n27502, n27545;
    
    LUT4 i3_3_lut_rep_352_4_lut (.A(count[12]), .B(n31576), .C(n29365), 
         .D(count[13]), .Z(n31495)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_352_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[0]), .B(n31578), .C(n31579), .D(n31577), 
         .Z(n29286)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX prev_in_46 (.D(n1170), .SP(n33386), .CK(debug_c_c), .Q(n1158));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i22476_3_lut_3_lut_4_lut (.A(n29110), .B(n31441), .C(n33381), 
         .D(n31439), .Z(n29402)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i22476_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i21_3_lut_rep_297_4_lut_4_lut (.A(n27607), .B(n31495), .C(count[9]), 
         .D(n10), .Z(n31440)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i21_3_lut_rep_297_4_lut_4_lut.init = 16'h1310;
    LUT4 i22010_3_lut_rep_465 (.A(n27607), .B(n31495), .C(count[9]), .Z(n33381)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i22010_3_lut_rep_465.init = 16'hecec;
    LUT4 i1_2_lut_rep_318_4_lut (.A(n31527), .B(count[13]), .C(n29365), 
         .D(count[9]), .Z(n31461)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_318_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(n10), .B(n33381), .C(n31461), .D(n28947), 
         .Z(n7)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31461), .C(n29286), 
         .D(n29110), .Z(n10_adj_204)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22012_3_lut_4_lut (.A(count[8]), .B(n31461), .C(n29110), .D(n29286), 
         .Z(n29568)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22012_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_rep_433 (.A(count[15]), .B(count[14]), .Z(n31576)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_433.init = 16'heeee;
    LUT4 i1_2_lut_rep_296_3_lut (.A(count[15]), .B(count[14]), .C(n27647), 
         .Z(n31439)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_296_3_lut.init = 16'hfefe;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_281 (.A(count[15]), .B(count[14]), .C(n5), 
         .D(n27647), .Z(n29403)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_281.init = 16'hfffe;
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    LUT4 i21957_2_lut_rep_384_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n31527)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i21957_2_lut_rep_384_3_lut.init = 16'hfefe;
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i14716_2_lut_rep_434 (.A(count[4]), .B(count[5]), .Z(n31577)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14716_2_lut_rep_434.init = 16'h8888;
    LUT4 i2_3_lut_rep_435 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n31578)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_435.init = 16'h8080;
    LUT4 i1_2_lut_rep_385_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n31528)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_385_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_436 (.A(count[6]), .B(count[7]), .Z(n31579)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_436.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), .Z(n29109)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_rep_383_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[5]), 
         .D(count[4]), .Z(n31526)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_rep_383_3_lut_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n33386), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1170));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(n1158), .B(n1170), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_298_3_lut (.A(count[9]), .B(n31495), .C(count[8]), 
         .Z(n31441)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_298_3_lut.init = 16'hfefe;
    CCU2D add_1774_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26502), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_17.INIT0 = 16'hd222;
    defparam add_1774_17.INIT1 = 16'h0000;
    defparam add_1774_17.INJECT1_0 = "NO";
    defparam add_1774_17.INJECT1_1 = "NO";
    CCU2D add_1774_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26501), 
          .COUT(n26502), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_15.INIT0 = 16'hd222;
    defparam add_1774_15.INIT1 = 16'hd222;
    defparam add_1774_15.INJECT1_0 = "NO";
    defparam add_1774_15.INJECT1_1 = "NO";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    CCU2D add_1774_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26500), 
          .COUT(n26501), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_13.INIT0 = 16'hd222;
    defparam add_1774_13.INIT1 = 16'hd222;
    defparam add_1774_13.INJECT1_0 = "NO";
    defparam add_1774_13.INJECT1_1 = "NO";
    LUT4 i22369_4_lut (.A(n31440), .B(n29523), .C(n28947), .D(n10_adj_204), 
         .Z(n29829)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22369_4_lut.init = 16'h3323;
    CCU2D add_1774_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26499), 
          .COUT(n26500), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_11.INIT0 = 16'hd222;
    defparam add_1774_11.INIT1 = 16'hd222;
    defparam add_1774_11.INJECT1_0 = "NO";
    defparam add_1774_11.INJECT1_1 = "NO";
    CCU2D add_1774_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26498), 
          .COUT(n26499), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_9.INIT0 = 16'hd222;
    defparam add_1774_9.INIT1 = 16'hd222;
    defparam add_1774_9.INJECT1_0 = "NO";
    defparam add_1774_9.INJECT1_1 = "NO";
    LUT4 i8_4_lut (.A(n31527), .B(n16), .C(count[13]), .D(count[11]), 
         .Z(n16912)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i8_4_lut.init = 16'h0004;
    LUT4 i7_4_lut (.A(count[10]), .B(n33385), .C(n26), .D(n29523), .Z(n16)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i7_4_lut.init = 16'h0040;
    CCU2D add_1774_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26497), 
          .COUT(n26498), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_7.INIT0 = 16'hd222;
    defparam add_1774_7.INIT1 = 16'hd222;
    defparam add_1774_7.INJECT1_0 = "NO";
    defparam add_1774_7.INJECT1_1 = "NO";
    LUT4 i33_3_lut (.A(n10), .B(n27607), .C(count[9]), .Z(n26)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_3_lut.init = 16'h3a3a;
    LUT4 i15395_2_lut (.A(n1092[7]), .B(n28947), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15395_2_lut.init = 16'h2222;
    CCU2D sub_73_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26754), 
          .S0(n1092[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_73_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_73_add_2_9.INIT1 = 16'h0000;
    defparam sub_73_add_2_9.INJECT1_0 = "NO";
    defparam sub_73_add_2_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n31461), .B(count[8]), .C(n31578), .D(n31526), 
         .Z(n28947)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(count[4]), .B(n31528), .C(count[8]), .D(n29109), 
         .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h8000;
    CCU2D sub_73_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26753), 
          .COUT(n26754), .S0(n1092[5]), .S1(n1092[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_73_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_73_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_73_add_2_7.INJECT1_0 = "NO";
    defparam sub_73_add_2_7.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_282 (.A(n27574), .B(n6), .C(count[8]), .D(n31577), 
         .Z(n27607)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_282.init = 16'hfefc;
    LUT4 i3_4_lut_adj_283 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27574)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_283.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_1774_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26496), 
          .COUT(n26497), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_5.INIT0 = 16'hd222;
    defparam add_1774_5.INIT1 = 16'hd222;
    defparam add_1774_5.INJECT1_0 = "NO";
    defparam add_1774_5.INJECT1_1 = "NO";
    CCU2D add_1774_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26495), 
          .COUT(n26496), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_3.INIT0 = 16'hd222;
    defparam add_1774_3.INIT1 = 16'hd222;
    defparam add_1774_3.INJECT1_0 = "NO";
    defparam add_1774_3.INJECT1_1 = "NO";
    CCU2D sub_73_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26752), 
          .COUT(n26753), .S0(n1092[3]), .S1(n1092[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_73_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_73_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_73_add_2_5.INJECT1_0 = "NO";
    defparam sub_73_add_2_5.INJECT1_1 = "NO";
    CCU2D add_1774_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29403), .B1(n1170), .C1(count[0]), .D1(n1158), .COUT(n26495), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_1.INIT0 = 16'hF000;
    defparam add_1774_1.INIT1 = 16'ha565;
    defparam add_1774_1.INJECT1_0 = "NO";
    defparam add_1774_1.INJECT1_1 = "NO";
    CCU2D sub_73_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26751), 
          .COUT(n26752), .S0(n1092[1]), .S1(n1092[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_73_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_73_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_73_add_2_3.INJECT1_0 = "NO";
    defparam sub_73_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_73_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26751), 
          .S1(n1092[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_73_add_2_1.INIT0 = 16'hF000;
    defparam sub_73_add_2_1.INIT1 = 16'h5555;
    defparam sub_73_add_2_1.INJECT1_0 = "NO";
    defparam sub_73_add_2_1.INJECT1_1 = "NO";
    LUT4 i21969_2_lut (.A(n1158), .B(n1170), .Z(n29523)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21969_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n29365)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_284 (.A(count[4]), .B(n29109), .C(count[3]), .D(n6_adj_205), 
         .Z(n29110)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_284.init = 16'hccc8;
    LUT4 i3300_2_lut (.A(count[1]), .B(count[2]), .Z(n6_adj_205)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3300_2_lut.init = 16'h8888;
    LUT4 i15394_2_lut (.A(n1092[6]), .B(n28947), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15394_2_lut.init = 16'h2222;
    LUT4 i15393_2_lut (.A(n1092[5]), .B(n28947), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15393_2_lut.init = 16'h2222;
    LUT4 i15392_2_lut (.A(n1092[4]), .B(n28947), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15392_2_lut.init = 16'h2222;
    LUT4 i15391_2_lut (.A(n1092[3]), .B(n28947), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15391_2_lut.init = 16'h2222;
    FD1P3AX valid_48 (.D(n29402), .SP(n27546), .CK(debug_c_c), .Q(n1164));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14513), .PD(n16912), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n29365), .D(n4), 
         .Z(n27647)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_285 (.A(n31579), .B(count[9]), .C(n27502), .D(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_285.init = 16'heccc;
    LUT4 i2_4_lut_adj_286 (.A(count[5]), .B(count[4]), .C(n6_adj_205), 
         .D(count[3]), .Z(n27502)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_286.init = 16'hfeee;
    LUT4 i15390_2_lut (.A(n1092[2]), .B(n28947), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15390_2_lut.init = 16'h2222;
    LUT4 i15389_2_lut (.A(n1092[1]), .B(n28947), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15389_2_lut.init = 16'h2222;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33386), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    LUT4 i22350_4_lut (.A(n31576), .B(n5), .C(n27647), .D(n27545), .Z(n29810)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22350_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_287 (.A(n33381), .B(n29523), .C(n7), .D(n29568), 
         .Z(n27545)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_287.init = 16'hdccc;
    LUT4 i15172_2_lut (.A(n1092[0]), .B(n28947), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15172_2_lut.init = 16'h2222;
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33386), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module SabertoothSerialPeripheral
//

module SabertoothSerialPeripheral (\read_size[0] , debug_c_c, n9378, n13907, 
            n31511, \databus[0] , \select[2] , read_value, n9541, 
            rw, n64, n31600, \register[0][7] , n31581, \reset_count[14] , 
            n22483, n11235, \databus[7] , \databus[6] , \databus[5] , 
            \databus[4] , \databus[3] , \databus[2] , \databus[1] , 
            \register_addr[0] , n31412, GND_net, n1155, n31536, \reset_count[8] , 
            \reset_count[7] , n29331, state, n29169, n31595, n31555, 
            n31575, n9, n33384, n31442, n31589, n35, n4180, \register_addr[5] , 
            n31463, n13916, \reset_count[11] , n21502, n27249, n29263, 
            n14782, n31529, n9296, n31462, motor_pwm_l_c, n8506, 
            n29785, select_clk, n2966, n107) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n9378;
    input n13907;
    input n31511;
    input \databus[0] ;
    input \select[2] ;
    output [7:0]read_value;
    input n9541;
    input rw;
    output n64;
    input n31600;
    output \register[0][7] ;
    output n31581;
    input \reset_count[14] ;
    input n22483;
    input n11235;
    input \databus[7] ;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    input \register_addr[0] ;
    input n31412;
    input GND_net;
    output n1155;
    input n31536;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29331;
    output [3:0]state;
    input n29169;
    input n31595;
    input n31555;
    input n31575;
    output n9;
    input n33384;
    input n31442;
    input n31589;
    input n35;
    output n4180;
    input \register_addr[5] ;
    input n31463;
    output n13916;
    input \reset_count[11] ;
    input n21502;
    input n27249;
    output n29263;
    input n14782;
    input n31529;
    output n9296;
    input n31462;
    output motor_pwm_l_c;
    output n8506;
    output n29785;
    output select_clk;
    input n2966;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n14966;
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire prev_select;
    wire [7:0]n28;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n29473, n9448;
    wire [31:0]n63;
    
    wire n31533, n27244, n9445;
    wire [7:0]n6204;
    
    FD1P3AX read_size__i1 (.D(n9378), .SP(n14966), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n13907), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam prev_select_138.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n28[0]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i16_2_lut (.A(\select[2] ), .B(rw), .Z(n64)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam i16_2_lut.init = 16'h8888;
    LUT4 i15387_4_lut_4_lut (.A(\register[1] [7]), .B(n31600), .C(n29473), 
         .D(n9448), .Z(n63[6])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i15387_4_lut_4_lut.init = 16'hffde;
    LUT4 i1_4_lut_4_lut (.A(\register[1] [7]), .B(n31600), .C(\register[1] [1]), 
         .D(n31533), .Z(n9448)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i1_4_lut_4_lut.init = 16'h2000;
    LUT4 i1_4_lut_4_lut_adj_280 (.A(\register[0][7] ), .B(n31600), .C(\register[0] [1]), 
         .D(n27244), .Z(n9445)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i1_4_lut_4_lut_adj_280.init = 16'h2000;
    LUT4 i1_2_lut_rep_438 (.A(\select[2] ), .B(prev_select), .Z(n31581)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_rep_438.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\select[2] ), .B(prev_select), .C(\reset_count[14] ), 
         .D(n22483), .Z(n14966)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    FD1P3IX register_0__i16 (.D(\databus[7] ), .SP(n11235), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n11235), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n11235), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n11235), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n11235), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n11235), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n11235), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n11235), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3IX register_0__i8 (.D(\databus[7] ), .SP(n13907), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[0][7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n13907), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n13907), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n13907), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n13907), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n13907), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n13907), .PD(n31511), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i2.GSR = "ENABLED";
    LUT4 mux_1915_Mux_7_i1_3_lut (.A(\register[0][7] ), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n6204[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1915_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n6204[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1915_Mux_5_i1_3_lut (.A(\register[0] [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n6204[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1915_Mux_4_i1_3_lut (.A(\register[0] [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n6204[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1915_Mux_3_i1_3_lut (.A(\register[0] [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n6204[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1915_Mux_2_i1_3_lut (.A(\register[0] [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n6204[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1915_Mux_1_i1_3_lut (.A(\register[0] [1]), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n6204[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_1_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i7 (.D(n6204[7]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6204[6]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6204[5]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6204[4]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6204[3]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n6204[2]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n6204[1]), .SP(n14966), .CD(n9541), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=528, LSE_RLINE=536 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1915_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n28[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1915_Mux_0_i1_3_lut.init = 16'hcaca;
    SabertoothSerial sserial (.debug_c_c(debug_c_c), .n31412(n31412), .GND_net(GND_net), 
            .\register[0][5] (\register[0] [5]), .n31600(n31600), .\register[0][6] (\register[0] [6]), 
            .\register[1][6] (\register[1] [6]), .n31533(n31533), .\register[1][7] (\register[1] [7]), 
            .\register[1][1] (\register[1] [1]), .\register[1][3] (\register[1] [3]), 
            .\register[1][5] (\register[1] [5]), .\register[1][4] (\register[1] [4]), 
            .\register[0][3] (\register[0] [3]), .\register[0][4] (\register[0] [4]), 
            .n1155(n1155), .n29473(n29473), .n89(n63[6]), .\register[0][7] (\register[0][7] ), 
            .n9445(n9445), .\register[1][2] (\register[1] [2]), .\register[0][2] (\register[0] [2]), 
            .n27244(n27244), .n31536(n31536), .n9448(n9448), .\register[0][1] (\register[0] [1]), 
            .\reset_count[8] (\reset_count[8] ), .\reset_count[7] (\reset_count[7] ), 
            .n29331(n29331), .state({state}), .n31511(n31511), .n29169(n29169), 
            .n31595(n31595), .n31555(n31555), .n31575(n31575), .n9(n9), 
            .n33384(n33384), .n31442(n31442), .n31589(n31589), .n35(n35), 
            .n4180(n4180), .rw(rw), .\register_addr[5] (\register_addr[5] ), 
            .n31463(n31463), .n13916(n13916), .\reset_count[11] (\reset_count[11] ), 
            .n21502(n21502), .n27249(n27249), .n29263(n29263), .n14782(n14782), 
            .n31529(n31529), .n9296(n9296), .n31462(n31462), .motor_pwm_l_c(motor_pwm_l_c), 
            .n22483(n22483), .\reset_count[14] (\reset_count[14] ), .n8506(n8506), 
            .n29785(n29785), .select_clk(select_clk), .n2966(n2966), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(142[19] 147[34])
    
endmodule
//
// Verilog Description of module SabertoothSerial
//

module SabertoothSerial (debug_c_c, n31412, GND_net, \register[0][5] , 
            n31600, \register[0][6] , \register[1][6] , n31533, \register[1][7] , 
            \register[1][1] , \register[1][3] , \register[1][5] , \register[1][4] , 
            \register[0][3] , \register[0][4] , n1155, n29473, n89, 
            \register[0][7] , n9445, \register[1][2] , \register[0][2] , 
            n27244, n31536, n9448, \register[0][1] , \reset_count[8] , 
            \reset_count[7] , n29331, state, n31511, n29169, n31595, 
            n31555, n31575, n9, n33384, n31442, n31589, n35, n4180, 
            rw, \register_addr[5] , n31463, n13916, \reset_count[11] , 
            n21502, n27249, n29263, n14782, n31529, n9296, n31462, 
            motor_pwm_l_c, n22483, \reset_count[14] , n8506, n29785, 
            select_clk, n2966, n107) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31412;
    input GND_net;
    input \register[0][5] ;
    input n31600;
    input \register[0][6] ;
    input \register[1][6] ;
    output n31533;
    input \register[1][7] ;
    input \register[1][1] ;
    input \register[1][3] ;
    input \register[1][5] ;
    input \register[1][4] ;
    input \register[0][3] ;
    input \register[0][4] ;
    output n1155;
    output n29473;
    input n89;
    input \register[0][7] ;
    input n9445;
    input \register[1][2] ;
    input \register[0][2] ;
    output n27244;
    input n31536;
    input n9448;
    input \register[0][1] ;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29331;
    output [3:0]state;
    input n31511;
    input n29169;
    input n31595;
    input n31555;
    input n31575;
    output n9;
    input n33384;
    input n31442;
    input n31589;
    input n35;
    output n4180;
    input rw;
    input \register_addr[5] ;
    input n31463;
    output n13916;
    input \reset_count[11] ;
    input n21502;
    input n27249;
    output n29263;
    input n14782;
    input n31529;
    output n9296;
    input n31462;
    output motor_pwm_l_c;
    input n22483;
    input \reset_count[14] ;
    output n8506;
    output n29785;
    output select_clk;
    input n2966;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [3:0]state_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    wire [3:0]n7808;
    wire [3:0]n16;
    
    wire n1, n31504, n10324;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(16[12:19])
    
    wire n14036, n31404, n29223, n20, n31586, n31471, n31588, 
        n31474, n12742, n31535, n31537, n12740, n28953, n6, n7, 
        n28310, n8;
    wire [7:0]n5504;
    wire [7:0]n5513;
    
    wire n12_adj_199;
    wire [31:0]n63;
    
    wire n6_adj_200, n11381, n11963, n12015, n12133, n24, n31502;
    
    FD1P3IX state__i1 (.D(n7808[1]), .SP(n31412), .CD(GND_net), .CK(debug_c_c), 
            .Q(state_c[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i1.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n16[0]), .CK(debug_c_c), .CD(GND_net), .Q(state_c[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 i3947_1_lut (.A(state_c[0]), .Z(n1)) /* synthesis lut_function=(!(A)) */ ;
    defparam i3947_1_lut.init = 16'h5555;
    LUT4 i15444_3_lut_4_lut (.A(\register[0][5] ), .B(n31504), .C(n31600), 
         .D(\register[0][6] ), .Z(n10324)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i15444_3_lut_4_lut.init = 16'hf8f0;
    FD1P3AX tx_data_i0_i0 (.D(n31404), .SP(n14036), .CK(debug_c_c), .Q(tx_data[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_390 (.A(\register[1][6] ), .B(n29223), .Z(n31533)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_390.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(\register[1][6] ), .B(n29223), .C(\register[1][7] ), 
         .D(\register[1][1] ), .Z(n20)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h80ff;
    LUT4 i5805_2_lut_rep_328_3_lut_4_lut (.A(\register[1][3] ), .B(n31586), 
         .C(\register[1][5] ), .D(\register[1][4] ), .Z(n31471)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5805_2_lut_rep_328_3_lut_4_lut.init = 16'h8000;
    LUT4 i5957_2_lut_rep_331_3_lut_4_lut (.A(\register[0][3] ), .B(n31588), 
         .C(\register[0][5] ), .D(\register[0][4] ), .Z(n31474)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5957_2_lut_rep_331_3_lut_4_lut.init = 16'h8000;
    LUT4 i5973_2_lut_3_lut_4_lut (.A(\register[0][3] ), .B(n31588), .C(\register[0][5] ), 
         .D(\register[0][4] ), .Z(n12742)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5973_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3IX send_31 (.D(n1), .SP(n31412), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1155));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam send_31.GSR = "ENABLED";
    LUT4 i4376_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n7808[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(34[6] 57[13])
    defparam i4376_2_lut.init = 16'h6666;
    LUT4 i21921_2_lut_3_lut_4_lut (.A(\register[1][4] ), .B(n31535), .C(\register[1][6] ), 
         .D(\register[1][5] ), .Z(n29473)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i21921_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i5971_2_lut_3_lut_4_lut (.A(\register[0][4] ), .B(n31537), .C(\register[0][6] ), 
         .D(\register[0][5] ), .Z(n12740)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5971_2_lut_3_lut_4_lut.init = 16'h78f0;
    PFUMX i30 (.BLUT(n28953), .ALUT(n6), .C0(n7), .Z(n28310));
    LUT4 i1_4_lut (.A(n31600), .B(\register[1][7] ), .C(n29473), .D(n8), 
         .Z(n28953)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut.init = 16'hffbf;
    LUT4 i1_2_lut (.A(\register[1][1] ), .B(n29223), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    PFUMX mux_1848_i7 (.BLUT(n89), .ALUT(n5504[6]), .C0(n7), .Z(n5513[6]));
    LUT4 i6_4_lut (.A(n31474), .B(n12_adj_199), .C(\register[0][7] ), 
         .D(state_c[1]), .Z(n6)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i6_4_lut.init = 16'h0080;
    PFUMX mux_1848_i2 (.BLUT(n63[1]), .ALUT(n5504[1]), .C0(n7), .Z(n5513[1]));
    LUT4 i5_4_lut (.A(\register[0][6] ), .B(state_c[0]), .C(n9445), .D(n31600), 
         .Z(n12_adj_199)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i5_4_lut.init = 16'h0002;
    PFUMX mux_1848_i3 (.BLUT(n63[2]), .ALUT(n5504[2]), .C0(n7), .Z(n5513[2]));
    LUT4 equal_16_i5_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(46[7:11])
    defparam equal_16_i5_2_lut.init = 16'hbbbb;
    LUT4 i3_4_lut (.A(\register[1][4] ), .B(\register[1][3] ), .C(\register[1][5] ), 
         .D(\register[1][2] ), .Z(n29223)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    PFUMX mux_1848_i4 (.BLUT(n63[3]), .ALUT(n5504[3]), .C0(n7), .Z(n5513[3]));
    LUT4 i4_4_lut (.A(\register[0][4] ), .B(\register[0][2] ), .C(\register[0][3] ), 
         .D(n6_adj_200), .Z(n27244)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_278 (.A(\register[0][5] ), .B(\register[0][6] ), .Z(n6_adj_200)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_278.init = 16'h8888;
    PFUMX mux_1848_i5 (.BLUT(n63[4]), .ALUT(n5504[4]), .C0(n7), .Z(n5513[4]));
    PFUMX mux_1848_i6 (.BLUT(n63[5]), .ALUT(n5504[5]), .C0(n7), .Z(n5513[5]));
    LUT4 i15046_4_lut (.A(n31536), .B(n11381), .C(n9445), .D(n10324), 
         .Z(n5504[6])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i15046_4_lut.init = 16'h3132;
    LUT4 i4391_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n11381)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i4391_2_lut.init = 16'heeee;
    LUT4 i15382_4_lut (.A(\register[1][2] ), .B(n9448), .C(n31600), .D(\register[1][1] ), 
         .Z(n63[1])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15382_4_lut.init = 16'hcdce;
    LUT4 i15038_4_lut (.A(n11963), .B(n11381), .C(n9445), .D(n31600), 
         .Z(n5504[1])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15038_4_lut.init = 16'h3032;
    LUT4 i5198_2_lut (.A(\register[0][2] ), .B(\register[0][1] ), .Z(n11963)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5198_2_lut.init = 16'h6666;
    LUT4 i15383_4_lut (.A(\register[1][3] ), .B(n9448), .C(n31600), .D(n31586), 
         .Z(n63[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15383_4_lut.init = 16'hcdce;
    LUT4 i15039_4_lut (.A(n12015), .B(n11381), .C(n9445), .D(n31600), 
         .Z(n5504[2])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15039_4_lut.init = 16'h3032;
    LUT4 i15384_4_lut (.A(\register[1][4] ), .B(n9448), .C(n31600), .D(n31535), 
         .Z(n63[3])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15384_4_lut.init = 16'hcdce;
    LUT4 i15040_4_lut (.A(n12133), .B(n11381), .C(n9445), .D(n31600), 
         .Z(n5504[3])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15040_4_lut.init = 16'h3032;
    LUT4 n20_bdd_4_lut (.A(n20), .B(n24), .C(n7), .D(n31600), .Z(n31404)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n20_bdd_4_lut.init = 16'h00ca;
    LUT4 i15385_4_lut (.A(\register[1][5] ), .B(n9448), .C(n31600), .D(n31502), 
         .Z(n63[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15385_4_lut.init = 16'hcdce;
    LUT4 i15041_4_lut (.A(n12742), .B(n11381), .C(n9445), .D(n31600), 
         .Z(n5504[4])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15041_4_lut.init = 16'h3032;
    LUT4 i15386_4_lut (.A(\register[1][6] ), .B(n9448), .C(n31600), .D(n31471), 
         .Z(n63[5])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15386_4_lut.init = 16'hcdce;
    LUT4 i4422_2_lut_rep_443 (.A(\register[1][2] ), .B(\register[1][1] ), 
         .Z(n31586)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4422_2_lut_rep_443.init = 16'h8888;
    LUT4 i5800_2_lut_rep_359_3_lut_4_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][4] ), .D(\register[1][3] ), .Z(n31502)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5800_2_lut_rep_359_3_lut_4_lut.init = 16'h8000;
    LUT4 i15043_4_lut (.A(n12740), .B(n11381), .C(n9445), .D(n31600), 
         .Z(n5504[5])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15043_4_lut.init = 16'h3032;
    LUT4 i4434_2_lut_rep_392_3_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][3] ), .Z(n31535)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i4434_2_lut_rep_392_3_lut.init = 16'h8080;
    LUT4 i5236_2_lut_rep_445 (.A(\register[0][2] ), .B(\register[0][1] ), 
         .Z(n31588)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5236_2_lut_rep_445.init = 16'h8888;
    LUT4 i5238_2_lut_rep_394_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n31537)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5238_2_lut_rep_394_3_lut.init = 16'h8080;
    LUT4 i5250_2_lut_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n12015)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i5250_2_lut_3_lut.init = 16'h7878;
    LUT4 i5955_2_lut_rep_361_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n31504)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5955_2_lut_rep_361_3_lut_4_lut.init = 16'h8000;
    LUT4 i5368_2_lut_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n12133)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5368_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3AX tx_data_i0_i1 (.D(n5513[1]), .SP(n14036), .CK(debug_c_c), 
            .Q(tx_data[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i2 (.D(n5513[2]), .SP(n14036), .CK(debug_c_c), 
            .Q(tx_data[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n5513[3]), .SP(n14036), .CK(debug_c_c), 
            .Q(tx_data[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n5513[4]), .SP(n14036), .CK(debug_c_c), 
            .Q(tx_data[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i5 (.D(n5513[5]), .SP(n14036), .CK(debug_c_c), 
            .Q(tx_data[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i6 (.D(n5513[6]), .SP(n14036), .CK(debug_c_c), 
            .Q(tx_data[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i7 (.D(n28310), .SP(n14036), .CK(debug_c_c), .Q(tx_data[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_279 (.A(n11381), .B(\register[0][1] ), .C(n27244), 
         .D(\register[0][7] ), .Z(n24)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;
    defparam i1_4_lut_adj_279.init = 16'h5111;
    \UARTTransmitter(baud_div=1250)  sender (.\reset_count[8] (\reset_count[8] ), 
            .\reset_count[7] (\reset_count[7] ), .n29331(n29331), .state({state}), 
            .n31511(n31511), .n29169(n29169), .n31595(n31595), .n31555(n31555), 
            .n31575(n31575), .n9(n9), .n33384(n33384), .n31442(n31442), 
            .n31589(n31589), .n35(n35), .n4180(n4180), .rw(rw), .\register_addr[5] (\register_addr[5] ), 
            .n31463(n31463), .n13916(n13916), .\reset_count[11] (\reset_count[11] ), 
            .n21502(n21502), .n27249(n27249), .n29263(n29263), .tx_data({tx_data}), 
            .n1155(n1155), .n14782(n14782), .n31529(n31529), .n9296(n9296), 
            .n31462(n31462), .motor_pwm_l_c(motor_pwm_l_c), .n22483(n22483), 
            .\reset_count[14] (\reset_count[14] ), .GND_net(GND_net), .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(63[26] 67[47])
    \ClockDividerP(factor=12000)  baud_gen (.GND_net(GND_net), .n8506(n8506), 
            .n29785(n29785), .n31511(n31511), .select_clk(select_clk), 
            .\state[0] (state_c[0]), .n14036(n14036), .n12(n16[0]), .debug_c_c(debug_c_c), 
            .n2966(n2966), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(21[25] 23[48])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=1250) 
//

module \UARTTransmitter(baud_div=1250)  (\reset_count[8] , \reset_count[7] , 
            n29331, state, n31511, n29169, n31595, n31555, n31575, 
            n9, n33384, n31442, n31589, n35, n4180, rw, \register_addr[5] , 
            n31463, n13916, \reset_count[11] , n21502, n27249, n29263, 
            tx_data, n1155, n14782, n31529, n9296, n31462, motor_pwm_l_c, 
            n22483, \reset_count[14] , GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29331;
    output [3:0]state;
    input n31511;
    input n29169;
    input n31595;
    input n31555;
    input n31575;
    output n9;
    input n33384;
    input n31442;
    input n31589;
    input n35;
    output n4180;
    input rw;
    input \register_addr[5] ;
    input n31463;
    output n13916;
    input \reset_count[11] ;
    input n21502;
    input n27249;
    output n29263;
    input [7:0]tx_data;
    input n1155;
    input n14782;
    input n31529;
    output n9296;
    input n31462;
    output motor_pwm_l_c;
    input n22483;
    input \reset_count[14] ;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n30718, n2780, n28470, n17, n30717, n30716;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9452, n7, n10, n104, n29770, n29771, n2, n29772, n29190, 
        n29191, n10_adj_198;
    
    LUT4 i1_2_lut (.A(\reset_count[8] ), .B(\reset_count[7] ), .Z(n29331)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX state__i0 (.D(n30718), .CK(bclk), .CD(n31511), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n31511), .B(state[3]), .C(state[2]), .D(n2780), 
         .Z(n28470)) /* synthesis lut_function=(!(A+(B (C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h1404;
    LUT4 i3_2_lut_4_lut (.A(n29169), .B(n31595), .C(n31555), .D(n31575), 
         .Z(n9)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i3_2_lut_4_lut.init = 16'h0200;
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 i2_3_lut_4_lut (.A(n33384), .B(n31442), .C(n31589), .D(n35), 
         .Z(n4180)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_4_lut_adj_274 (.A(rw), .B(n31442), .C(\register_addr[5] ), 
         .D(n31463), .Z(n13916)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_274.init = 16'h0004;
    PFUMX i22645 (.BLUT(n30717), .ALUT(n30716), .C0(state[2]), .Z(n30718));
    LUT4 i1_4_lut_adj_275 (.A(\reset_count[11] ), .B(n21502), .C(\reset_count[8] ), 
         .D(n27249), .Z(n29263)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_275.init = 16'h8880;
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9452), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;
    LUT4 state_1__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n30716)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(n1155), .Z(n30717)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8f0e;
    LUT4 i22210_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n29770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22210_3_lut.init = 16'hcaca;
    LUT4 i22211_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n29771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22211_3_lut.init = 16'hcaca;
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n29772), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15421_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15421_4_lut.init = 16'hfcee;
    FD1P3AX state__i3 (.D(n28470), .SP(n14782), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(n31511), .B(state[2]), .C(state[3]), .D(n2780), 
         .Z(n29190)) /* synthesis lut_function=(!(A+(B (C+(D))+!B !(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1104;
    LUT4 i4_4_lut (.A(n31442), .B(n31529), .C(n31589), .D(rw), .Z(n9296)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i4_4_lut.init = 16'h0008;
    FD1P3AX state__i2 (.D(n29190), .SP(n14782), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n29191), .SP(n14782), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(state[1]), .B(n31462), .C(state[0]), .Z(n29191)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n31511), .CK(bclk), .Q(motor_pwm_l_c)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    PFUMX i22212 (.BLUT(n29770), .ALUT(n29771), .C0(state[1]), .Z(n29772));
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9452), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9452), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9452), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9452), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9452), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9452), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9452), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_276 (.A(state[1]), .B(state[0]), .Z(n2780)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_276.init = 16'h8888;
    LUT4 i5_4_lut (.A(state[3]), .B(n10_adj_198), .C(n22483), .D(state[1]), 
         .Z(n9452)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i5_4_lut.init = 16'h0040;
    LUT4 i4_4_lut_adj_277 (.A(\reset_count[14] ), .B(state[2]), .C(state[0]), 
         .D(n1155), .Z(n10_adj_198)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i4_4_lut_adj_277.init = 16'h0200;
    \ClockDividerP(factor=1250)  baud_gen (.GND_net(GND_net), .bclk(bclk), 
            .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=1250) 
//

module \ClockDividerP(factor=1250)  (GND_net, bclk, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output bclk;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27144;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n8541, n27143, n27142, n27141, n27140, n27139, n27138, 
        n27137, n27136, n27135, n27134, n27133, n27132, n27131, 
        n27130, n27066;
    wire [31:0]n102;
    
    wire n27065, n29843, n45, n52, n46, n16804, n50, n42, n27064, 
        n27063, n27062, n27061, n48, n38, n27060, n27059, n27058, 
        n44, n30, n29621, n27057, n27056, n27055, n27054, n27053, 
        n27052, n27051;
    
    CCU2D add_19625_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27144), 
          .S1(n8541));
    defparam add_19625_32.INIT0 = 16'h5555;
    defparam add_19625_32.INIT1 = 16'h0000;
    defparam add_19625_32.INJECT1_0 = "NO";
    defparam add_19625_32.INJECT1_1 = "NO";
    CCU2D add_19625_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27143), .COUT(n27144));
    defparam add_19625_30.INIT0 = 16'h5555;
    defparam add_19625_30.INIT1 = 16'h5555;
    defparam add_19625_30.INJECT1_0 = "NO";
    defparam add_19625_30.INJECT1_1 = "NO";
    CCU2D add_19625_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27142), .COUT(n27143));
    defparam add_19625_28.INIT0 = 16'h5555;
    defparam add_19625_28.INIT1 = 16'h5555;
    defparam add_19625_28.INJECT1_0 = "NO";
    defparam add_19625_28.INJECT1_1 = "NO";
    CCU2D add_19625_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27141), .COUT(n27142));
    defparam add_19625_26.INIT0 = 16'h5555;
    defparam add_19625_26.INIT1 = 16'h5555;
    defparam add_19625_26.INJECT1_0 = "NO";
    defparam add_19625_26.INJECT1_1 = "NO";
    CCU2D add_19625_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27140), .COUT(n27141));
    defparam add_19625_24.INIT0 = 16'h5555;
    defparam add_19625_24.INIT1 = 16'h5555;
    defparam add_19625_24.INJECT1_0 = "NO";
    defparam add_19625_24.INJECT1_1 = "NO";
    CCU2D add_19625_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27139), .COUT(n27140));
    defparam add_19625_22.INIT0 = 16'h5555;
    defparam add_19625_22.INIT1 = 16'h5555;
    defparam add_19625_22.INJECT1_0 = "NO";
    defparam add_19625_22.INJECT1_1 = "NO";
    CCU2D add_19625_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27138), .COUT(n27139));
    defparam add_19625_20.INIT0 = 16'h5555;
    defparam add_19625_20.INIT1 = 16'h5555;
    defparam add_19625_20.INJECT1_0 = "NO";
    defparam add_19625_20.INJECT1_1 = "NO";
    CCU2D add_19625_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27137), .COUT(n27138));
    defparam add_19625_18.INIT0 = 16'h5555;
    defparam add_19625_18.INIT1 = 16'h5555;
    defparam add_19625_18.INJECT1_0 = "NO";
    defparam add_19625_18.INJECT1_1 = "NO";
    CCU2D add_19625_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27136), .COUT(n27137));
    defparam add_19625_16.INIT0 = 16'h5555;
    defparam add_19625_16.INIT1 = 16'h5555;
    defparam add_19625_16.INJECT1_0 = "NO";
    defparam add_19625_16.INJECT1_1 = "NO";
    CCU2D add_19625_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27135), .COUT(n27136));
    defparam add_19625_14.INIT0 = 16'h5555;
    defparam add_19625_14.INIT1 = 16'h5555;
    defparam add_19625_14.INJECT1_0 = "NO";
    defparam add_19625_14.INJECT1_1 = "NO";
    CCU2D add_19625_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27134), .COUT(n27135));
    defparam add_19625_12.INIT0 = 16'h5555;
    defparam add_19625_12.INIT1 = 16'h5555;
    defparam add_19625_12.INJECT1_0 = "NO";
    defparam add_19625_12.INJECT1_1 = "NO";
    CCU2D add_19625_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27133), .COUT(n27134));
    defparam add_19625_10.INIT0 = 16'h5aaa;
    defparam add_19625_10.INIT1 = 16'h5555;
    defparam add_19625_10.INJECT1_0 = "NO";
    defparam add_19625_10.INJECT1_1 = "NO";
    CCU2D add_19625_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27132), 
          .COUT(n27133));
    defparam add_19625_8.INIT0 = 16'h5555;
    defparam add_19625_8.INIT1 = 16'h5555;
    defparam add_19625_8.INJECT1_0 = "NO";
    defparam add_19625_8.INJECT1_1 = "NO";
    CCU2D add_19625_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27131), 
          .COUT(n27132));
    defparam add_19625_6.INIT0 = 16'h5aaa;
    defparam add_19625_6.INIT1 = 16'h5aaa;
    defparam add_19625_6.INJECT1_0 = "NO";
    defparam add_19625_6.INJECT1_1 = "NO";
    CCU2D add_19625_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27130), 
          .COUT(n27131));
    defparam add_19625_4.INIT0 = 16'h5555;
    defparam add_19625_4.INIT1 = 16'h5aaa;
    defparam add_19625_4.INJECT1_0 = "NO";
    defparam add_19625_4.INJECT1_1 = "NO";
    CCU2D add_19625_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27130));
    defparam add_19625_2.INIT0 = 16'h1000;
    defparam add_19625_2.INIT1 = 16'h5555;
    defparam add_19625_2.INJECT1_0 = "NO";
    defparam add_19625_2.INJECT1_1 = "NO";
    FD1S3AX clk_o_14 (.D(n8541), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2680_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27066), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_33.INIT1 = 16'h0000;
    defparam count_2680_add_4_33.INJECT1_0 = "NO";
    defparam count_2680_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27065), .COUT(n27066), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_31.INJECT1_0 = "NO";
    defparam count_2680_add_4_31.INJECT1_1 = "NO";
    LUT4 i22385_4_lut (.A(n29843), .B(n45), .C(n52), .D(n46), .Z(n16804)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22385_4_lut.init = 16'h0002;
    LUT4 i22383_4_lut (.A(count[13]), .B(n50), .C(n42), .D(count[3]), 
         .Z(n29843)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22383_4_lut.init = 16'h0001;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n45)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    CCU2D count_2680_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27064), .COUT(n27065), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_29.INJECT1_0 = "NO";
    defparam count_2680_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27063), .COUT(n27064), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_27.INJECT1_0 = "NO";
    defparam count_2680_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27062), .COUT(n27063), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_25.INJECT1_0 = "NO";
    defparam count_2680_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27061), .COUT(n27062), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_23.INJECT1_0 = "NO";
    defparam count_2680_add_4_23.INJECT1_1 = "NO";
    LUT4 i24_4_lut (.A(count[30]), .B(n48), .C(n38), .D(count[14]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(count[24]), .B(count[4]), .C(count[1]), .D(count[27]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i18_4_lut.init = 16'hfffe;
    CCU2D count_2680_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27060), .COUT(n27061), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_21.INJECT1_0 = "NO";
    defparam count_2680_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27059), .COUT(n27060), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_19.INJECT1_0 = "NO";
    defparam count_2680_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27058), .COUT(n27059), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_17.INJECT1_0 = "NO";
    defparam count_2680_add_4_17.INJECT1_1 = "NO";
    LUT4 i22_4_lut (.A(count[28]), .B(n44), .C(n30), .D(count[18]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(count[31]), .B(count[5]), .C(n29621), .D(count[6]), 
         .Z(n42)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i14_4_lut.init = 16'hbfff;
    CCU2D count_2680_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27057), .COUT(n27058), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_15.INJECT1_0 = "NO";
    defparam count_2680_add_4_15.INJECT1_1 = "NO";
    LUT4 i16_4_lut (.A(count[16]), .B(count[21]), .C(count[11]), .D(count[25]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[2]), .B(count[8]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(count[20]), .B(count[23]), .C(count[15]), .D(count[29]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20_4_lut.init = 16'hfffe;
    CCU2D count_2680_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27056), .COUT(n27057), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_13.INJECT1_0 = "NO";
    defparam count_2680_add_4_13.INJECT1_1 = "NO";
    LUT4 i10_2_lut (.A(count[19]), .B(count[22]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i22062_3_lut (.A(count[10]), .B(count[0]), .C(count[7]), .Z(n29621)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22062_3_lut.init = 16'h8080;
    CCU2D count_2680_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27055), .COUT(n27056), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_11.INJECT1_0 = "NO";
    defparam count_2680_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27054), .COUT(n27055), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_9.INJECT1_0 = "NO";
    defparam count_2680_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27053), .COUT(n27054), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_7.INJECT1_0 = "NO";
    defparam count_2680_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27052), .COUT(n27053), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_5.INJECT1_0 = "NO";
    defparam count_2680_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27051), .COUT(n27052), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_3.INJECT1_0 = "NO";
    defparam count_2680_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27051), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_1.INIT0 = 16'hF000;
    defparam count_2680_add_4_1.INIT1 = 16'h0555;
    defparam count_2680_add_4_1.INJECT1_0 = "NO";
    defparam count_2680_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2680__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i0.GSR = "ENABLED";
    FD1S3IX count_2680__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i1.GSR = "ENABLED";
    FD1S3IX count_2680__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i2.GSR = "ENABLED";
    FD1S3IX count_2680__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i3.GSR = "ENABLED";
    FD1S3IX count_2680__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i4.GSR = "ENABLED";
    FD1S3IX count_2680__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i5.GSR = "ENABLED";
    FD1S3IX count_2680__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i6.GSR = "ENABLED";
    FD1S3IX count_2680__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i7.GSR = "ENABLED";
    FD1S3IX count_2680__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i8.GSR = "ENABLED";
    FD1S3IX count_2680__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i9.GSR = "ENABLED";
    FD1S3IX count_2680__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i10.GSR = "ENABLED";
    FD1S3IX count_2680__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i11.GSR = "ENABLED";
    FD1S3IX count_2680__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i12.GSR = "ENABLED";
    FD1S3IX count_2680__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i13.GSR = "ENABLED";
    FD1S3IX count_2680__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i14.GSR = "ENABLED";
    FD1S3IX count_2680__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i15.GSR = "ENABLED";
    FD1S3IX count_2680__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i16.GSR = "ENABLED";
    FD1S3IX count_2680__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i17.GSR = "ENABLED";
    FD1S3IX count_2680__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i18.GSR = "ENABLED";
    FD1S3IX count_2680__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i19.GSR = "ENABLED";
    FD1S3IX count_2680__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i20.GSR = "ENABLED";
    FD1S3IX count_2680__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i21.GSR = "ENABLED";
    FD1S3IX count_2680__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i22.GSR = "ENABLED";
    FD1S3IX count_2680__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i23.GSR = "ENABLED";
    FD1S3IX count_2680__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i24.GSR = "ENABLED";
    FD1S3IX count_2680__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i25.GSR = "ENABLED";
    FD1S3IX count_2680__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i26.GSR = "ENABLED";
    FD1S3IX count_2680__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i27.GSR = "ENABLED";
    FD1S3IX count_2680__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i28.GSR = "ENABLED";
    FD1S3IX count_2680__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i29.GSR = "ENABLED";
    FD1S3IX count_2680__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i30.GSR = "ENABLED";
    FD1S3IX count_2680__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000) 
//

module \ClockDividerP(factor=12000)  (GND_net, n8506, n29785, n31511, 
            select_clk, \state[0] , n14036, n12, debug_c_c, n2966, 
            n107) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n8506;
    output n29785;
    input n31511;
    output select_clk;
    input \state[0] ;
    output n14036;
    output n12;
    input debug_c_c;
    input n2966;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27157;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27156, n27155, n27154, n27153, n27152, n27151, n27150, 
        n27149, n27148, n27147, n27146, n27145, n27781, n15, n20, 
        n16, n27, n40, n36, n28, n18, n38, n32;
    wire [31:0]n134;
    
    wire n34, n24, n27050, n27049, n27048, n27047, n27046, n27045, 
        n27044, n27043, n27042, n27041, n27040, n27039, n27038, 
        n27037, n27036, n27035;
    
    CCU2D add_19624_28 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27157), 
          .S1(n8506));
    defparam add_19624_28.INIT0 = 16'h5555;
    defparam add_19624_28.INIT1 = 16'h0000;
    defparam add_19624_28.INJECT1_0 = "NO";
    defparam add_19624_28.INJECT1_1 = "NO";
    CCU2D add_19624_26 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27156), .COUT(n27157));
    defparam add_19624_26.INIT0 = 16'h5555;
    defparam add_19624_26.INIT1 = 16'h5555;
    defparam add_19624_26.INJECT1_0 = "NO";
    defparam add_19624_26.INJECT1_1 = "NO";
    CCU2D add_19624_24 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27155), .COUT(n27156));
    defparam add_19624_24.INIT0 = 16'h5555;
    defparam add_19624_24.INIT1 = 16'h5555;
    defparam add_19624_24.INJECT1_0 = "NO";
    defparam add_19624_24.INJECT1_1 = "NO";
    CCU2D add_19624_22 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27154), .COUT(n27155));
    defparam add_19624_22.INIT0 = 16'h5555;
    defparam add_19624_22.INIT1 = 16'h5555;
    defparam add_19624_22.INJECT1_0 = "NO";
    defparam add_19624_22.INJECT1_1 = "NO";
    CCU2D add_19624_20 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27153), .COUT(n27154));
    defparam add_19624_20.INIT0 = 16'h5555;
    defparam add_19624_20.INIT1 = 16'h5555;
    defparam add_19624_20.INJECT1_0 = "NO";
    defparam add_19624_20.INJECT1_1 = "NO";
    CCU2D add_19624_18 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27152), .COUT(n27153));
    defparam add_19624_18.INIT0 = 16'h5555;
    defparam add_19624_18.INIT1 = 16'h5555;
    defparam add_19624_18.INJECT1_0 = "NO";
    defparam add_19624_18.INJECT1_1 = "NO";
    CCU2D add_19624_16 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27151), .COUT(n27152));
    defparam add_19624_16.INIT0 = 16'h5555;
    defparam add_19624_16.INIT1 = 16'h5555;
    defparam add_19624_16.INJECT1_0 = "NO";
    defparam add_19624_16.INJECT1_1 = "NO";
    CCU2D add_19624_14 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27150), .COUT(n27151));
    defparam add_19624_14.INIT0 = 16'h5555;
    defparam add_19624_14.INIT1 = 16'h5555;
    defparam add_19624_14.INJECT1_0 = "NO";
    defparam add_19624_14.INJECT1_1 = "NO";
    CCU2D add_19624_12 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27149), .COUT(n27150));
    defparam add_19624_12.INIT0 = 16'h5555;
    defparam add_19624_12.INIT1 = 16'h5555;
    defparam add_19624_12.INJECT1_0 = "NO";
    defparam add_19624_12.INJECT1_1 = "NO";
    CCU2D add_19624_10 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27148), .COUT(n27149));
    defparam add_19624_10.INIT0 = 16'h5555;
    defparam add_19624_10.INIT1 = 16'h5555;
    defparam add_19624_10.INJECT1_0 = "NO";
    defparam add_19624_10.INJECT1_1 = "NO";
    CCU2D add_19624_8 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27147), .COUT(n27148));
    defparam add_19624_8.INIT0 = 16'h5555;
    defparam add_19624_8.INIT1 = 16'h5aaa;
    defparam add_19624_8.INJECT1_0 = "NO";
    defparam add_19624_8.INJECT1_1 = "NO";
    CCU2D add_19624_6 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27146), .COUT(n27147));
    defparam add_19624_6.INIT0 = 16'h5aaa;
    defparam add_19624_6.INIT1 = 16'h5aaa;
    defparam add_19624_6.INJECT1_0 = "NO";
    defparam add_19624_6.INJECT1_1 = "NO";
    CCU2D add_19624_4 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27145), 
          .COUT(n27146));
    defparam add_19624_4.INIT0 = 16'h5555;
    defparam add_19624_4.INIT1 = 16'h5aaa;
    defparam add_19624_4.INJECT1_0 = "NO";
    defparam add_19624_4.INJECT1_1 = "NO";
    CCU2D add_19624_2 (.A0(count[5]), .B0(count[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27145));
    defparam add_19624_2.INIT0 = 16'h7000;
    defparam add_19624_2.INIT1 = 16'h5aaa;
    defparam add_19624_2.INJECT1_0 = "NO";
    defparam add_19624_2.INJECT1_1 = "NO";
    LUT4 i22325_4_lut (.A(n27781), .B(n15), .C(n20), .D(n16), .Z(n29785)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i22325_4_lut.init = 16'h4000;
    LUT4 i20_4_lut (.A(n27), .B(n40), .C(n36), .D(n28), .Z(n27781)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[11]), .B(count[10]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(count[9]), .B(n18), .C(count[6]), .D(count[7]), 
         .Z(n20)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(count[1]), .B(count[4]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i22356_2_lut_4_lut (.A(n31511), .B(select_clk), .C(n8506), .D(\state[0] ), 
         .Z(n14036)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i22356_2_lut_4_lut.init = 16'h0010;
    LUT4 i5968_2_lut_4_lut (.A(n31511), .B(select_clk), .C(n8506), .D(\state[0] ), 
         .Z(n12)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i5968_2_lut_4_lut.init = 16'hef10;
    LUT4 i6_2_lut (.A(count[28]), .B(count[12]), .Z(n27)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[5]), .B(n38), .C(n32), .D(count[20]), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(count[8]), .B(count[25]), .C(count[15]), .D(count[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_4_lut.init = 16'hfffe;
    FD1S3IX count_2679__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2966), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i0.GSR = "ENABLED";
    LUT4 i7_2_lut (.A(count[17]), .B(count[24]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i7_4_lut (.A(count[13]), .B(count[2]), .C(count[3]), .D(count[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i17_4_lut (.A(count[29]), .B(n34), .C(n24), .D(count[14]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(count[22]), .B(count[21]), .C(count[31]), .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(count[16]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[19]), .B(count[18]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    FD1S3AX clk_o_14 (.D(n107), .CK(debug_c_c), .Q(select_clk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=25, LSE_RCOL=48, LSE_LLINE=21, LSE_RLINE=23 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2679_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27050), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_33.INIT1 = 16'h0000;
    defparam count_2679_add_4_33.INJECT1_0 = "NO";
    defparam count_2679_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27049), .COUT(n27050), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_31.INJECT1_0 = "NO";
    defparam count_2679_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27048), .COUT(n27049), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_29.INJECT1_0 = "NO";
    defparam count_2679_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27047), .COUT(n27048), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_27.INJECT1_0 = "NO";
    defparam count_2679_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27046), .COUT(n27047), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_25.INJECT1_0 = "NO";
    defparam count_2679_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27045), .COUT(n27046), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_23.INJECT1_0 = "NO";
    defparam count_2679_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27044), .COUT(n27045), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_21.INJECT1_0 = "NO";
    defparam count_2679_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27043), .COUT(n27044), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_19.INJECT1_0 = "NO";
    defparam count_2679_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27042), .COUT(n27043), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_17.INJECT1_0 = "NO";
    defparam count_2679_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27041), .COUT(n27042), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_15.INJECT1_0 = "NO";
    defparam count_2679_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27040), .COUT(n27041), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_13.INJECT1_0 = "NO";
    defparam count_2679_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27039), .COUT(n27040), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_11.INJECT1_0 = "NO";
    defparam count_2679_add_4_11.INJECT1_1 = "NO";
    FD1S3IX count_2679__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2966), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i1.GSR = "ENABLED";
    CCU2D count_2679_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27038), .COUT(n27039), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_9.INJECT1_0 = "NO";
    defparam count_2679_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27037), .COUT(n27038), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_7.INJECT1_0 = "NO";
    defparam count_2679_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27036), .COUT(n27037), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_5.INJECT1_0 = "NO";
    defparam count_2679_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27035), .COUT(n27036), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_3.INJECT1_0 = "NO";
    defparam count_2679_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27035), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_1.INIT0 = 16'hF000;
    defparam count_2679_add_4_1.INIT1 = 16'h0555;
    defparam count_2679_add_4_1.INJECT1_0 = "NO";
    defparam count_2679_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2679__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2966), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i2.GSR = "ENABLED";
    FD1S3IX count_2679__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2966), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i3.GSR = "ENABLED";
    FD1S3IX count_2679__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2966), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i4.GSR = "ENABLED";
    FD1S3IX count_2679__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2966), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i5.GSR = "ENABLED";
    FD1S3IX count_2679__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2966), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i6.GSR = "ENABLED";
    FD1S3IX count_2679__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2966), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i7.GSR = "ENABLED";
    FD1S3IX count_2679__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2966), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i8.GSR = "ENABLED";
    FD1S3IX count_2679__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2966), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i9.GSR = "ENABLED";
    FD1S3IX count_2679__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i10.GSR = "ENABLED";
    FD1S3IX count_2679__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i11.GSR = "ENABLED";
    FD1S3IX count_2679__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i12.GSR = "ENABLED";
    FD1S3IX count_2679__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i13.GSR = "ENABLED";
    FD1S3IX count_2679__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i14.GSR = "ENABLED";
    FD1S3IX count_2679__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i15.GSR = "ENABLED";
    FD1S3IX count_2679__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i16.GSR = "ENABLED";
    FD1S3IX count_2679__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i17.GSR = "ENABLED";
    FD1S3IX count_2679__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i18.GSR = "ENABLED";
    FD1S3IX count_2679__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i19.GSR = "ENABLED";
    FD1S3IX count_2679__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i20.GSR = "ENABLED";
    FD1S3IX count_2679__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i21.GSR = "ENABLED";
    FD1S3IX count_2679__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i22.GSR = "ENABLED";
    FD1S3IX count_2679__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i23.GSR = "ENABLED";
    FD1S3IX count_2679__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i24.GSR = "ENABLED";
    FD1S3IX count_2679__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i25.GSR = "ENABLED";
    FD1S3IX count_2679__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i26.GSR = "ENABLED";
    FD1S3IX count_2679__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i27.GSR = "ENABLED";
    FD1S3IX count_2679__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i28.GSR = "ENABLED";
    FD1S3IX count_2679__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i29.GSR = "ENABLED";
    FD1S3IX count_2679__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i30.GSR = "ENABLED";
    FD1S3IX count_2679__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2966), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (register_addr, debug_c_c, databus, 
            \select[7] , n33389, \select[5] , \select[4] , \select[3] , 
            \select[2] , \select[1] , databus_out, n13833, \sendcount[1] , 
            n31555, n29300, n31532, n29199, debug_c_5, n31496, rw, 
            n31425, prev_select, n31427, n31595, n31469, n31465, 
            n31426, \register[1][19] , n59, n31500, \register[1][20] , 
            n57, \register[1][26] , n45, force_pause, \register[2] , 
            \register[1][0] , n97, n31503, prev_select_adj_5, n31511, 
            n13940, n1491, n29169, n29294, n29068, n29292, n31435, 
            n303, n56, n29293, n29065, n29055, n29052, n29064, 
            n29062, n29049, n224, n3921, n29051, n29053, n27751, 
            n29066, n29056, n29067, n29070, n29071, n27752, n29069, 
            n29057, n29058, n29063, n29059, n29257, n29061, n29054, 
            n29050, n29048, n29060, n29047, prev_select_adj_6, n2846, 
            n66, \register[0][2] , read_value, n33384, n2, n31464, 
            n2_adj_7, n2_adj_8, n2_adj_9, n2_adj_10, n31540, n31449, 
            n31477, n31470, n2_adj_11, n2_adj_12, n2_adj_13, n31473, 
            n2_adj_14, n2_adj_15, n2_adj_16, n2_adj_17, n2_adj_18, 
            n2_adj_19, n2_adj_20, n2_adj_21, n2_adj_22, n2_adj_23, 
            n3, n3_adj_24, n3_adj_25, n31589, n31476, n3_adj_26, 
            n3_adj_27, n3_adj_28, n3_adj_29, n3_adj_30, n2_adj_31, 
            n2_adj_32, n2_adj_33, n2_adj_34, n2_adj_35, n2_adj_36, 
            n31482, n14453, n9537, n35, n27464, n33383, n31445, 
            debug_c_7, \read_size[2] , n29234, n31444, n52, n31442, 
            n29236, n176, n31448, n31570, n16012, n31456, n31581, 
            n13907, n11235, n31434, n30305, n29220, n31525, n31419, 
            n30303, \control_reg[7] , n1, n31529, n31539, n13155, 
            n13, n18, n14, \reg_size[2] , n31587, n31590, n27441, 
            \control_reg[7]_adj_37 , n31600, n32, n4, n5833, prev_select_adj_38, 
            \reset_count[14] , n22483, n2869, n224_adj_91, n4094, 
            n31575, \read_value[7]_adj_71 , n2_adj_72, \read_value[5]_adj_73 , 
            n2_adj_74, n31472, \read_value[4]_adj_75 , n2_adj_76, \read_value[6]_adj_77 , 
            n2_adj_78, \read_value[3]_adj_79 , n2_adj_80, \read_value[2]_adj_81 , 
            n2_adj_82, \read_value[0]_adj_83 , n2_adj_84, n27444, n34, 
            n29256, n9330, n1485, \register[0][5] , expansion5_c, 
            \register[1][5] , debug_c_2, n1488, debug_c_3, n9378, 
            n29491, prev_select_adj_85, \steps_reg[7] , n11, debug_c_4, 
            n31501, n6005, \steps_reg[5] , n14_adj_86, \register[0][4] , 
            expansion4_out, \register[1][4] , timeout_pause, \steps_reg[6] , 
            n13_adj_87, \register[0][7] , n31536, clk_1Hz, signal_light_c, 
            \steps_reg[3] , n12, \control_reg[4] , \div_factor_reg[4] , 
            \steps_reg[4] , \control_reg[7]_adj_88 , n8635, n13947, 
            n12368, n9300, n14522, n4006, n31406, n27679, n27483, 
            n32_adj_89, n16764, n9, n9304, prev_select_adj_90, n16763, 
            n6002, n27427, n28826, n8653, \state[3] , \state[1] , 
            \state[0] , n1155, n73, \reset_count[7] , \reset_count[6] , 
            \reset_count[5] , n27249, n11072, GND_net, uart_rx_c) /* synthesis syn_module_defined=1 */ ;
    output [7:0]register_addr;
    input debug_c_c;
    input [31:0]databus;
    output \select[7] ;
    input n33389;
    output \select[5] ;
    output \select[4] ;
    output \select[3] ;
    output \select[2] ;
    output \select[1] ;
    output [31:0]databus_out;
    input n13833;
    output \sendcount[1] ;
    output n31555;
    output n29300;
    output n31532;
    output n29199;
    output debug_c_5;
    output n31496;
    output rw;
    output n31425;
    input prev_select;
    output n31427;
    output n31595;
    output n31469;
    output n31465;
    output n31426;
    input \register[1][19] ;
    output n59;
    input n31500;
    input \register[1][20] ;
    output n57;
    input \register[1][26] ;
    output n45;
    input force_pause;
    input [31:0]\register[2] ;
    input \register[1][0] ;
    output n97;
    output n31503;
    input prev_select_adj_5;
    input n31511;
    output n13940;
    output n1491;
    input n29169;
    output n29294;
    output n29068;
    output n29292;
    output n31435;
    output n303;
    output n56;
    output n29293;
    output n29065;
    output n29055;
    output n29052;
    output n29064;
    output n29062;
    output n29049;
    input [31:0]n224;
    output [31:0]n3921;
    output n29051;
    output n29053;
    output n27751;
    output n29066;
    output n29056;
    output n29067;
    output n29070;
    output n29071;
    output n27752;
    output n29069;
    output n29057;
    output n29058;
    output n29063;
    output n29059;
    output n29257;
    output n29061;
    output n29054;
    output n29050;
    output n29048;
    output n29060;
    output n29047;
    input prev_select_adj_6;
    output n2846;
    output n66;
    input \register[0][2] ;
    input [31:0]read_value;
    output n33384;
    output n2;
    output n31464;
    output n2_adj_7;
    output n2_adj_8;
    output n2_adj_9;
    output n2_adj_10;
    input n31540;
    output n31449;
    output n31477;
    output n31470;
    output n2_adj_11;
    output n2_adj_12;
    output n2_adj_13;
    output n31473;
    output n2_adj_14;
    output n2_adj_15;
    output n2_adj_16;
    output n2_adj_17;
    output n2_adj_18;
    output n2_adj_19;
    output n2_adj_20;
    output n2_adj_21;
    output n2_adj_22;
    output n2_adj_23;
    output n3;
    output n3_adj_24;
    output n3_adj_25;
    output n31589;
    output n31476;
    output n3_adj_26;
    output n3_adj_27;
    output n3_adj_28;
    output n3_adj_29;
    output n3_adj_30;
    output n2_adj_31;
    output n2_adj_32;
    output n2_adj_33;
    output n2_adj_34;
    output n2_adj_35;
    output n2_adj_36;
    output n31482;
    input n14453;
    output n9537;
    input n35;
    input n27464;
    input n33383;
    output n31445;
    output debug_c_7;
    input \read_size[2] ;
    output n29234;
    output n31444;
    output n52;
    output n31442;
    input n29236;
    output n176;
    output n31448;
    output n31570;
    output n16012;
    output n31456;
    input n31581;
    output n13907;
    output n11235;
    output n31434;
    output n30305;
    output n29220;
    output n31525;
    output n31419;
    output n30303;
    input \control_reg[7] ;
    output n1;
    output n31529;
    output n31539;
    input n13155;
    input n13;
    input n18;
    input n14;
    input \reg_size[2] ;
    input n31587;
    input n31590;
    input n27441;
    input \control_reg[7]_adj_37 ;
    output n31600;
    output n32;
    output n4;
    output n5833;
    input prev_select_adj_38;
    input \reset_count[14] ;
    input n22483;
    output n2869;
    input [31:0]n224_adj_91;
    output [31:0]n4094;
    output n31575;
    input \read_value[7]_adj_71 ;
    output n2_adj_72;
    input \read_value[5]_adj_73 ;
    output n2_adj_74;
    input n31472;
    input \read_value[4]_adj_75 ;
    output n2_adj_76;
    input \read_value[6]_adj_77 ;
    output n2_adj_78;
    input \read_value[3]_adj_79 ;
    output n2_adj_80;
    input \read_value[2]_adj_81 ;
    output n2_adj_82;
    input \read_value[0]_adj_83 ;
    output n2_adj_84;
    input n27444;
    output n34;
    output n29256;
    output n9330;
    output n1485;
    input \register[0][5] ;
    input expansion5_c;
    input \register[1][5] ;
    output debug_c_2;
    output n1488;
    output debug_c_3;
    output n9378;
    output n29491;
    input prev_select_adj_85;
    input \steps_reg[7] ;
    output n11;
    output debug_c_4;
    output n31501;
    output n6005;
    input \steps_reg[5] ;
    output n14_adj_86;
    input \register[0][4] ;
    input expansion4_out;
    input \register[1][4] ;
    input timeout_pause;
    input \steps_reg[6] ;
    output n13_adj_87;
    input \register[0][7] ;
    output n31536;
    input clk_1Hz;
    output signal_light_c;
    input \steps_reg[3] ;
    output n12;
    input \control_reg[4] ;
    input \div_factor_reg[4] ;
    input \steps_reg[4] ;
    input \control_reg[7]_adj_88 ;
    output n8635;
    output n13947;
    output n12368;
    output n9300;
    output n14522;
    output n4006;
    output n31406;
    output n27679;
    input n27483;
    output n32_adj_89;
    output n16764;
    input n9;
    output n9304;
    input prev_select_adj_90;
    output n16763;
    output n6002;
    output n27427;
    output n28826;
    output n8653;
    input \state[3] ;
    input \state[1] ;
    input \state[0] ;
    input n1155;
    output n73;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n27249;
    output n11072;
    input GND_net;
    input uart_rx_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire n33383 /* synthesis nomerge= */ ;
    
    wire n2805;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [31:0]n1473;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n29357, n5, n5_adj_39, n29021, n27597, n5_adj_40, n29022, 
        n27538;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n31475;
    wire [4:0]n15;
    
    wire n15667, n5_adj_41, n29023, n27548, n31400, n31399, n31646, 
        n16685, n31643, n2807;
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    wire [7:0]n5824;
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n31610, n33380, n15679;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n31468;
    wire [7:0]n2215;
    
    wire n15782, n30707, n5_adj_42, n29024, n27556;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n9471, n28592, n31447, n30823, n5_adj_43, n29027, n27524, 
        n31612, n31611, n31543, n31548, n10, n31553, n11_c, n11_adj_44, 
        n11_adj_45, n11_adj_46, n11_adj_47, n11_adj_48, n11_adj_49, 
        n11_adj_50, n31618, n31617, n31949, n31951, n2746, n16769, 
        n31621, n31620, n31624, n31623, n30302, n28916, n29389, 
        n31627, n31626, n31630, n31629, n15674, n1926, n31633, 
        n31632, n31645, n15670;
    wire [4:0]n17;
    
    wire n27681, n31636, n31635, n27433, n31639, n31638, n31608, 
        n31609, n31641, n31644, n9_adj_53, n31583, n31505, n31642, 
        n31423, n5_adj_54, n29025, n27504, n31450, n31541;
    wire [3:0]n1869;
    
    wire n31414, n31422, n31585, n31534, n4_c, n31622;
    wire [7:0]n9241;
    
    wire n4_adj_55, n31625, n29358, n4_adj_56, n31613, n4_adj_57, 
        n31631, n13489, n29204, n31486, n5_adj_58, n29028, n27472, 
        n31453, n14_c, n5_adj_59, n29031, n27532, n29018, n29255, 
        n29019, n29020, n5_adj_60, n29030, n27557, n31507, escape, 
        n10974, n30304, n5_adj_62, n29026, n27491, n4_adj_63, n31637, 
        n4_adj_64, n31634, n5_adj_65, n29032, n27555, n5_adj_69, 
        n29033, n27554, n2224, n29034, n29029, n5_adj_71, n27551, 
        n29035, n29036, n31544, n5_adj_77, n27550, n29360, n29037, 
        n31584, n31640, n30705, n30706, n5_adj_82, n27500, n7, 
        n30339, n29573, n38, n4_adj_85, n31628, n29038, n29039, 
        n29040, n29041, n29042, n29043, n29044, n5_adj_88, n27543, 
        n5_adj_89, n27533, n29045, n30822, n5_adj_95, n27426, n29014, 
        n5_adj_97, n27478, n29017, n29015, n5_adj_98, n27610, n29016, 
        n31552, n27625, n5_adj_102, n27496, n5_adj_103, n27513, 
        n29361, n5_adj_107, n27512, n31599, n57_adj_109, n31478, 
        n5_adj_110, n27476, n11_adj_111, n11_adj_112, n11_adj_113, 
        n11_adj_114, n5_adj_115, n27511, n31551, n11_adj_116, n11_adj_117, 
        n11_adj_118, n11_adj_119, n5_adj_120, n27510, send, n5_adj_121, 
        n27465, n31512, n1874, n31549, n31550, n9_adj_122, n5_adj_123, 
        n27505, n6, n5_adj_124, n27499, n31514, n7_adj_125, n31522, 
        n28666, n28658, n31538, n28616, n31523, n29276, n28, n29230, 
        n28614, n28618, n28620, n28662, n15678, n1_adj_126, n6_adj_127, 
        n28612, n28660, n15781, n31506, n28624, n28608, n28610, 
        n30340, n28586, n28622, n28606, n5_adj_130, n27601, n5_adj_131, 
        n27599, n15666, n16684, n27602, n31415, n13788, n31580, 
        n30341, n30733, n13_adj_151, busy, n11202, n19331;
    wire [7:0]register_addr_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    
    wire n12349, n79, n159, n8, n10_adj_157, n13041, n45_adj_163, 
        n112, n28899, n25, n19, n12_adj_172, n6_adj_173, n29162, 
        n28692, n16767, n13464, n12481, n29228, n1578, n1584, 
        n1585, n11216, n12347, n28604, n8_adj_182, n8_adj_185, n7_adj_186, 
        n29647, n29559, n29423, n30735;
    
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    LUT4 select_2129_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1473[4]), 
         .C(rx_data[2]), .D(n29357), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut (.A(databus[3]), .B(n5_adj_39), .C(n1473[13]), .D(n29021), 
         .Z(n27597)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 select_2129_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1473[4]), 
         .C(rx_data[3]), .D(n29357), .Z(n5_adj_39)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_82 (.A(databus[4]), .B(n5_adj_40), .C(n1473[13]), 
         .D(n29022), .Z(n27538)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_82.init = 16'hffec;
    LUT4 select_2129_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1473[4]), 
         .C(rx_data[4]), .D(n29357), .Z(n5_adj_40)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_20_i5_4_lut.init = 16'h88c0;
    FD1P3AX sendcount__i0 (.D(n15[0]), .SP(n31475), .CK(debug_c_c), .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    FD1S3IX select__i7 (.D(n15667), .CK(debug_c_c), .CD(n33389), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_83 (.A(databus[5]), .B(n5_adj_41), .C(n1473[13]), 
         .D(n29023), .Z(n27548)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_83.init = 16'hffec;
    FD1S3IX select__i5 (.D(n31400), .CK(debug_c_c), .CD(n33389), .Q(\select[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i5.GSR = "ENABLED";
    FD1S3IX select__i4 (.D(n31399), .CK(debug_c_c), .CD(n33389), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1S3IX select__i3 (.D(n31646), .CK(debug_c_c), .CD(n33389), .Q(\select[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i3.GSR = "ENABLED";
    FD1S3IX select__i2 (.D(n16685), .CK(debug_c_c), .CD(n33389), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1S3IX select__i1 (.D(n31643), .CK(debug_c_c), .CD(n33389), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    LUT4 select_2129_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1473[4]), 
         .C(rx_data[5]), .D(n29357), .Z(n5_adj_41)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_21_i5_4_lut.init = 16'h88c0;
    FD1P3AX esc_data_i0_i4 (.D(n5824[4]), .SP(n13833), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n5824[2]), .SP(n13833), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n5824[1]), .SP(n13833), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    FD1S3IX bufcount__i3 (.D(n31610), .CK(debug_c_c), .CD(n33389), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n33380), .CK(debug_c_c), .CD(n33389), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n15679), .CK(debug_c_c), .CD(n33389), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2215[4]), .SP(n31468), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2215[3]), .SP(n31468), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2215[1]), .SP(n31468), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n2215[0]), .SP(n31468), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n15782), .CK(debug_c_c), .CD(n33389), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n30707), .SP(n13833), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2807), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_84 (.A(databus[6]), .B(n5_adj_42), .C(n1473[13]), 
         .D(n29024), .Z(n27556)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_84.init = 16'hffec;
    FD1P3IX buffer_0___i1 (.D(n28592), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 select_2129_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1473[4]), 
         .C(rx_data[6]), .D(n29357), .Z(n5_adj_42)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_22_i5_4_lut.init = 16'h88c0;
    FD1P3IX sendcount__i4 (.D(n30823), .SP(n31475), .CD(n31447), .CK(debug_c_c), 
            .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_85 (.A(databus[7]), .B(n5_adj_43), .C(n1473[13]), 
         .D(n29027), .Z(n27524)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_85.init = 16'hffec;
    LUT4 i22191_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n31612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22191_then_3_lut.init = 16'hcaca;
    LUT4 i22191_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n31611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22191_else_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(register_addr[1]), .B(n31555), .C(register_addr[4]), 
         .D(n31543), .Z(n29300)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut.init = 16'h0002;
    LUT4 i2_2_lut_3_lut_4_lut (.A(register_addr[1]), .B(n31555), .C(n31532), 
         .D(register_addr[4]), .Z(n29199)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i5_3_lut_4_lut (.A(n31548), .B(n1473[12]), .C(n10), .D(n1473[9]), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_3_lut_4_lut.init = 16'hfffe;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n31553), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_c)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_86 (.A(bufcount[0]), .B(n31553), .C(rx_data[1]), 
         .D(\buffer[0] [1]), .Z(n11_adj_44)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_86.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_87 (.A(bufcount[0]), .B(n31553), .C(rx_data[2]), 
         .D(\buffer[0] [2]), .Z(n11_adj_45)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_87.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_88 (.A(bufcount[0]), .B(n31553), .C(\buffer[0] [3]), 
         .D(rx_data[3]), .Z(n11_adj_46)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_88.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_89 (.A(bufcount[0]), .B(n31553), .C(\buffer[0] [4]), 
         .D(rx_data[4]), .Z(n11_adj_47)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_89.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_90 (.A(bufcount[0]), .B(n31553), .C(\buffer[0] [5]), 
         .D(rx_data[5]), .Z(n11_adj_48)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_90.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_91 (.A(bufcount[0]), .B(n31553), .C(\buffer[0] [6]), 
         .D(rx_data[6]), .Z(n11_adj_49)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_91.init = 16'hf1e0;
    LUT4 i20_2_lut_rep_282_3_lut_4_lut (.A(\select[4] ), .B(n31496), .C(rw), 
         .D(register_addr[5]), .Z(n31425)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i20_2_lut_rep_282_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_284_3_lut_4_lut (.A(\select[4] ), .B(n31496), .C(prev_select), 
         .D(register_addr[5]), .Z(n31427)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_284_3_lut_4_lut.init = 16'h0800;
    LUT4 i24_3_lut_4_lut_adj_92 (.A(bufcount[0]), .B(n31553), .C(rx_data[7]), 
         .D(\buffer[0] [7]), .Z(n11_adj_50)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_92.init = 16'hfe10;
    LUT4 i1_2_lut_rep_326_3_lut_4_lut (.A(register_addr[4]), .B(n31595), 
         .C(register_addr[5]), .D(n31555), .Z(n31469)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_rep_326_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(\sendcount[1] ), .C(sendcount[0]), 
         .D(sendcount[2]), .Z(n31618)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_rep_322_3_lut_4_lut (.A(register_addr[4]), .B(n31595), 
         .C(\select[4] ), .D(n31555), .Z(n31465)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_rep_322_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(\sendcount[1] ), .C(sendcount[0]), 
         .D(sendcount[2]), .Z(n31617)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 n31949_bdd_4_lut (.A(n31949), .B(n1473[4]), .C(n31951), .D(bufcount[2]), 
         .Z(n33380)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n31949_bdd_4_lut.init = 16'heef0;
    LUT4 i1_2_lut_3_lut (.A(register_addr[0]), .B(n31426), .C(\register[1][19] ), 
         .Z(n59)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i15752_3_lut_rep_325 (.A(n2746), .B(n31500), .C(n1473[18]), .Z(n31468)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15752_3_lut_rep_325.init = 16'hc8c8;
    LUT4 i22346_2_lut_3_lut (.A(n2746), .B(n31500), .C(n1473[18]), .Z(n16769)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i22346_2_lut_3_lut.init = 16'h0808;
    LUT4 i22176_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n31621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22176_then_3_lut.init = 16'hcaca;
    LUT4 i22176_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n31620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22176_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_93 (.A(register_addr[0]), .B(n31426), .C(\register[1][20] ), 
         .Z(n57)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_93.init = 16'h2020;
    LUT4 i22179_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n31624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22179_then_3_lut.init = 16'hcaca;
    LUT4 i22179_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n31623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22179_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_94 (.A(register_addr[0]), .B(n31426), .C(\register[1][26] ), 
         .Z(n45)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_94.init = 16'h2020;
    LUT4 force_pause_bdd_4_lut (.A(force_pause), .B(register_addr[0]), .C(register_addr[1]), 
         .D(\register[2] [1]), .Z(n30302)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam force_pause_bdd_4_lut.init = 16'h3e0e;
    LUT4 i1_2_lut_3_lut_adj_95 (.A(register_addr[0]), .B(n31426), .C(\register[1][0] ), 
         .Z(n97)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_95.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_96 (.A(\buffer[0] [1]), .B(n28916), .C(\buffer[0] [2]), 
         .Z(n29389)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i1_2_lut_3_lut_adj_96.init = 16'hefef;
    LUT4 i22194_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n31627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22194_then_3_lut.init = 16'hcaca;
    LUT4 i22194_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n31626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22194_else_3_lut.init = 16'hcaca;
    LUT4 i22197_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n31630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22197_then_3_lut.init = 16'hcaca;
    LUT4 i22197_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n31629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22197_else_3_lut.init = 16'hcaca;
    LUT4 \buffer_0[[0__bdd_4_lut_22978  (.A(\buffer[0] [0]), .B(n29389), 
         .C(n15674), .D(n1926), .Z(n31399)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam \buffer_0[[0__bdd_4_lut_22978 .init = 16'h11f0;
    LUT4 i22200_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n31633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22200_then_3_lut.init = 16'hcaca;
    LUT4 i22200_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n31632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22200_else_3_lut.init = 16'hcaca;
    LUT4 n13750_bdd_4_lut_then_3_lut_4_lut (.A(\buffer[0] [2]), .B(\buffer[0] [0]), 
         .C(n28916), .D(\buffer[0] [1]), .Z(n31645)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam n13750_bdd_4_lut_then_3_lut_4_lut.init = 16'h0400;
    LUT4 \buffer_0[[0__bdd_4_lut  (.A(\buffer[0] [0]), .B(n29389), .C(n15670), 
         .D(n1926), .Z(n31400)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam \buffer_0[[0__bdd_4_lut .init = 16'h22f0;
    FD1P3IX sendcount__i3 (.D(n17[3]), .SP(n31475), .CD(n31447), .CK(debug_c_c), 
            .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3IX sendcount__i2 (.D(n17[2]), .SP(n31475), .CD(n31447), .CK(debug_c_c), 
            .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n17[1]), .SP(n31475), .CD(n31447), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 i22424_3_lut_4_lut (.A(\buffer[0] [1]), .B(n28916), .C(\buffer[0] [0]), 
         .D(\buffer[0] [2]), .Z(n27681)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i22424_3_lut_4_lut.init = 16'h2000;
    LUT4 i22203_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n31636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22203_then_3_lut.init = 16'hcaca;
    LUT4 i22203_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n31635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22203_else_3_lut.init = 16'hcaca;
    LUT4 i22464_3_lut_4_lut (.A(\buffer[0] [1]), .B(n28916), .C(\buffer[0] [0]), 
         .D(\buffer[0] [2]), .Z(n27433)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i22464_3_lut_4_lut.init = 16'h0002;
    LUT4 i22639_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n31639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22639_then_3_lut.init = 16'hcaca;
    LUT4 i22639_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n31638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22639_else_3_lut.init = 16'hcaca;
    LUT4 i8897_else_4_lut (.A(bufcount[3]), .B(n1473[0]), .C(n1473[3]), 
         .D(n1473[4]), .Z(n31608)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8897_else_4_lut.init = 16'h0002;
    LUT4 i8897_then_4_lut (.A(bufcount[3]), .B(n1473[0]), .C(n1473[3]), 
         .D(n1473[4]), .Z(n31609)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8897_then_4_lut.init = 16'haaa2;
    LUT4 n13673_bdd_4_lut_else_3_lut (.A(\select[1] ), .B(n1473[8]), .C(n1473[0]), 
         .Z(n31641)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam n13673_bdd_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(\select[4] ), .B(n31503), .C(prev_select_adj_5), 
         .D(n31511), .Z(n13940)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 n13750_bdd_4_lut_else_3_lut (.A(\select[3] ), .B(n1473[8]), .C(n1473[0]), 
         .Z(n31644)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam n13750_bdd_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i15750_3_lut_rep_332 (.A(n1473[13]), .B(n31500), .C(n1491), .Z(n31475)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15750_3_lut_rep_332.init = 16'hc8c8;
    LUT4 i14816_4_lut (.A(sendcount[3]), .B(n9_adj_53), .C(sendcount[2]), 
         .D(n31583), .Z(n17[3])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(271[10:37])
    defparam i14816_4_lut.init = 16'h4888;
    LUT4 i22349_2_lut_rep_304_3_lut (.A(n1473[13]), .B(n31500), .C(n1491), 
         .Z(n31447)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i22349_2_lut_rep_304_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(n31505), .C(\register[2] [31]), 
         .D(n29169), .Z(n29294)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_97 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [28]), .D(n29169), .Z(n29068)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_97.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_98 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [29]), .D(n29169), .Z(n29292)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_98.init = 16'h1000;
    LUT4 select_2129_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1473[4]), 
         .C(rx_data[7]), .D(n29357), .Z(n5_adj_43)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 n13673_bdd_4_lut_then_3_lut_4_lut (.A(\buffer[0] [2]), .B(\buffer[0] [0]), 
         .C(n28916), .D(\buffer[0] [1]), .Z(n31642)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam n13673_bdd_4_lut_then_3_lut_4_lut.init = 16'h0004;
    LUT4 register_addr_1__bdd_3_lut_22611_rep_292_4_lut (.A(register_addr[2]), 
         .B(n31505), .C(register_addr[0]), .D(register_addr[1]), .Z(n31435)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam register_addr_1__bdd_3_lut_22611_rep_292_4_lut.init = 16'h0110;
    LUT4 i21971_2_lut_rep_280_3_lut_4_lut (.A(register_addr[2]), .B(n31505), 
         .C(rw), .D(register_addr[1]), .Z(n31423)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i21971_2_lut_rep_280_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_99 (.A(register_addr[2]), .B(n31505), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n303)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_99.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_100 (.A(register_addr[2]), .B(n31505), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_100.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_101 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [30]), .D(n29169), .Z(n29293)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_101.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_102 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [4]), .D(n29169), .Z(n29065)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_102.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_103 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [5]), .D(n29169), .Z(n29055)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_103.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_104 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [6]), .D(n29169), .Z(n29052)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_104.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_105 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [7]), .D(n29169), .Z(n29064)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_105.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_106 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [8]), .D(n29169), .Z(n29062)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_106.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_107 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [9]), .D(n29169), .Z(n29049)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_107.init = 16'h1000;
    LUT4 i2_4_lut_adj_108 (.A(databus[8]), .B(n5_adj_54), .C(n1473[13]), 
         .D(n29025), .Z(n27504)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_108.init = 16'hffec;
    LUT4 i3351_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n31450), .C(n31541), 
         .D(bufcount[0]), .Z(n1869[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3351_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    LUT4 mux_1553_i13_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[12]), 
         .D(n224[12]), .Z(n3921[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_109 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [10]), .D(n29169), .Z(n29051)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_109.init = 16'h1000;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n31585), .B(n31534), .C(n4_c), 
         .D(n31622), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n31585), .B(n31534), .C(n4_adj_55), 
         .D(n31625), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 select_2129_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1473[4]), 
         .C(rx_data[0]), .D(n29358), .Z(n5_adj_54)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n31585), .B(n31534), .C(n4_adj_56), 
         .D(n31613), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n31585), .B(n31534), .C(n4_adj_57), 
         .D(n31631), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_4_lut_adj_110 (.A(n31553), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n13489), .Z(n29204)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_110.init = 16'h0e00;
    LUT4 i22113_2_lut_rep_343_4_lut (.A(register_addr[5]), .B(n31595), .C(register_addr[4]), 
         .D(n31555), .Z(n31486)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22113_2_lut_rep_343_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_111 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [11]), .D(n29169), .Z(n29053)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_111.init = 16'h1000;
    LUT4 i22341_3_lut_4_lut (.A(n31555), .B(register_addr[1]), .C(register_addr[4]), 
         .D(n31532), .Z(n27751)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i22341_3_lut_4_lut.init = 16'h0010;
    LUT4 i2_4_lut_adj_112 (.A(databus[9]), .B(n5_adj_58), .C(n1473[13]), 
         .D(n29028), .Z(n27472)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_112.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_113 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [12]), .D(n29169), .Z(n29066)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_113.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_114 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [13]), .D(n29169), .Z(n29056)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_114.init = 16'h1000;
    LUT4 select_2129_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1473[4]), 
         .C(rx_data[1]), .D(n29358), .Z(n5_adj_58)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_115 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [14]), .D(n29169), .Z(n29067)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_115.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_116 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [15]), .D(n29169), .Z(n29070)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_116.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_117 (.A(n1473[3]), .B(n31453), .C(n1473[13]), 
         .Z(n14_c)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_117.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_118 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [16]), .D(n29169), .Z(n29071)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_118.init = 16'h1000;
    LUT4 i22338_3_lut_4_lut (.A(n31555), .B(register_addr[1]), .C(register_addr[4]), 
         .D(n31543), .Z(n27752)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i22338_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_119 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [17]), .D(n29169), .Z(n29069)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_119.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_120 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [18]), .D(n29169), .Z(n29057)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_120.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_121 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [19]), .D(n29169), .Z(n29058)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_121.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_122 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [20]), .D(n29169), .Z(n29063)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_122.init = 16'h1000;
    LUT4 i2_4_lut_adj_123 (.A(databus[10]), .B(n5_adj_59), .C(n1473[13]), 
         .D(n29031), .Z(n27532)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_123.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_124 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [21]), .D(n29169), .Z(n29059)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_124.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_125 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [0]), 
         .Z(n29018)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_125.init = 16'h8080;
    LUT4 select_2129_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1473[4]), 
         .C(rx_data[2]), .D(n29358), .Z(n5_adj_59)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i1_3_lut_4_lut (.A(n31555), .B(register_addr[1]), .C(n29255), 
         .D(n31595), .Z(n29257)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_126 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [22]), .D(n29169), .Z(n29061)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_126.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_127 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [1]), 
         .Z(n29019)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_127.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_128 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [23]), .D(n29169), .Z(n29054)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_128.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_129 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [24]), .D(n29169), .Z(n29050)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_129.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_130 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [2]), 
         .Z(n29020)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_130.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_131 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [3]), 
         .Z(n29021)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_131.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_132 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [25]), .D(n29169), .Z(n29048)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_132.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_133 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [26]), .D(n29169), .Z(n29060)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_133.init = 16'h1000;
    FD1P3AX rw_498 (.D(n1473[10]), .SP(n2805), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_134 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [4]), 
         .Z(n29022)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_134.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_135 (.A(register_addr[2]), .B(n31505), 
         .C(\register[2] [27]), .D(n29169), .Z(n29047)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_135.init = 16'h1000;
    LUT4 i2_4_lut_adj_136 (.A(databus[11]), .B(n5_adj_60), .C(n1473[13]), 
         .D(n29030), .Z(n27557)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_136.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_adj_137 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [5]), 
         .Z(n29023)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_137.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_138 (.A(n31507), .B(prev_select_adj_6), 
         .C(\select[4] ), .D(n31511), .Z(n2846)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_138.init = 16'h0010;
    LUT4 i1_2_lut (.A(\select[5] ), .B(rw), .Z(n66)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(454[7:9])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_139 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [6]), 
         .Z(n29024)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_139.init = 16'h8080;
    FD1S3AX escape_501 (.D(n10974), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_140 (.A(n1473[3]), .B(n31453), .C(\buffer[2] [7]), 
         .Z(n29027)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_140.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_141 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [0]), 
         .Z(n29025)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_141.init = 16'h8080;
    LUT4 select_2129_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1473[4]), 
         .C(rx_data[3]), .D(n29358), .Z(n5_adj_60)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_142 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [1]), 
         .Z(n29028)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_142.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_143 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [2]), 
         .Z(n29031)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_143.init = 16'h8080;
    LUT4 \register_0[[2__bdd_4_lut  (.A(\register[0][2] ), .B(register_addr[0]), 
         .C(register_addr[1]), .D(\register[2] [2]), .Z(n30304)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam \register_0[[2__bdd_4_lut .init = 16'h3e0e;
    LUT4 i2_4_lut_adj_144 (.A(databus[12]), .B(n5_adj_62), .C(n1473[13]), 
         .D(n29026), .Z(n27491)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_144.init = 16'hffec;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n31585), .B(n31534), .C(n4_adj_63), 
         .D(n31637), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 select_2129_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1473[4]), 
         .C(rx_data[4]), .D(n29358), .Z(n5_adj_62)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n31585), .B(n31534), .C(n4_adj_64), 
         .D(n31634), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_adj_145 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [3]), 
         .Z(n29030)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_145.init = 16'h8080;
    LUT4 Select_4243_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[23]), .D(n33384), .Z(n2)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4243_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_146 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [4]), 
         .Z(n29026)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_146.init = 16'h8080;
    LUT4 i2_4_lut_adj_147 (.A(databus[13]), .B(n5_adj_65), .C(n1473[13]), 
         .D(n29032), .Z(n27555)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_147.init = 16'hffec;
    LUT4 select_2129_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1473[4]), 
         .C(rx_data[5]), .D(n29358), .Z(n5_adj_65)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 i14702_2_lut_rep_321_3_lut_4_lut (.A(register_addr[5]), .B(n31595), 
         .C(\select[3] ), .D(register_addr[4]), .Z(n31464)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i14702_2_lut_rep_321_3_lut_4_lut.init = 16'he0f0;
    LUT4 Select_4246_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[22]), .D(n33384), .Z(n2_adj_7)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4246_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4249_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[21]), .D(n33384), .Z(n2_adj_8)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4249_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4252_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[20]), .D(n33384), .Z(n2_adj_9)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4252_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_148 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [5]), 
         .Z(n29032)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_148.init = 16'h8080;
    LUT4 i2_4_lut_adj_149 (.A(databus[14]), .B(n5_adj_69), .C(n1473[13]), 
         .D(n29033), .Z(n27554)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_149.init = 16'hffec;
    LUT4 Select_4237_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[25]), .D(rw), .Z(n2_adj_10)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4237_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i22_1_lut_rep_306_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31595), 
         .C(n31540), .D(register_addr[4]), .Z(n31449)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i22_1_lut_rep_306_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_adj_150 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [6]), 
         .Z(n29033)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_150.init = 16'h8080;
    LUT4 i1_2_lut_adj_151 (.A(n1473[16]), .B(n1473[19]), .Z(n2224)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_151.init = 16'heeee;
    LUT4 select_2129_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1473[4]), 
         .C(rx_data[6]), .D(n29358), .Z(n5_adj_69)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_152 (.A(n1473[3]), .B(n31453), .C(\buffer[3] [7]), 
         .Z(n29034)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_152.init = 16'h8080;
    LUT4 i1_2_lut_rep_334_3_lut_4_lut (.A(register_addr[5]), .B(n31595), 
         .C(n31540), .D(register_addr[4]), .Z(n31477)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_334_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_153 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [0]), 
         .Z(n29029)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_153.init = 16'h8080;
    LUT4 i2_4_lut_adj_154 (.A(databus[15]), .B(n5_adj_71), .C(n1473[13]), 
         .D(n29034), .Z(n27551)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_154.init = 16'hffec;
    LUT4 i15036_2_lut_rep_327_3_lut_4_lut (.A(register_addr[5]), .B(n31595), 
         .C(\select[3] ), .D(register_addr[4]), .Z(n31470)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i15036_2_lut_rep_327_3_lut_4_lut.init = 16'h1000;
    LUT4 select_2129_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1473[4]), 
         .C(rx_data[7]), .D(n29358), .Z(n5_adj_71)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4240_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[24]), .D(n33384), .Z(n2_adj_11)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4240_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4255_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[19]), .D(n33384), .Z(n2_adj_12)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4255_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_155 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [1]), 
         .Z(n29035)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_155.init = 16'h8080;
    LUT4 Select_4258_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[18]), .D(rw), .Z(n2_adj_13)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4258_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_156 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [2]), 
         .Z(n29036)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_156.init = 16'h8080;
    LUT4 i1_2_lut_rep_330_3_lut_4_lut (.A(register_addr[5]), .B(n31595), 
         .C(\select[4] ), .D(n31544), .Z(n31473)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_330_3_lut_4_lut.init = 16'h0010;
    LUT4 Select_4261_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[17]), .D(rw), .Z(n2_adj_14)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4261_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4264_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[16]), .D(rw), .Z(n2_adj_15)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4264_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_157 (.A(databus[16]), .B(n5_adj_77), .C(n1473[13]), 
         .D(n29029), .Z(n27550)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_157.init = 16'hffec;
    LUT4 select_2129_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1473[4]), 
         .C(rx_data[0]), .D(n29360), .Z(n5_adj_77)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4267_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[15]), .D(rw), .Z(n2_adj_16)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4267_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4270_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[14]), .D(rw), .Z(n2_adj_17)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4270_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_158 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [3]), 
         .Z(n29037)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_158.init = 16'h8080;
    LUT4 Select_4273_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[13]), .D(rw), .Z(n2_adj_18)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4273_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 n30705_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n31584), .C(n31640), 
         .D(n30705), .Z(n30706)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n30705_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 Select_4276_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[12]), .D(rw), .Z(n2_adj_19)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4276_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_159 (.A(databus[17]), .B(n5_adj_82), .C(n1473[13]), 
         .D(n29035), .Z(n27500)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_159.init = 16'hffec;
    LUT4 select_2129_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1473[4]), 
         .C(rx_data[1]), .D(n29360), .Z(n5_adj_82)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut (.A(n1473[15]), .B(n7), .C(n30339), .D(n29573), .Z(n38)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'haaa8;
    LUT4 Select_4279_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[11]), .D(rw), .Z(n2_adj_20)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4279_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4282_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[10]), .D(rw), .Z(n2_adj_21)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4282_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n31585), .B(n31534), .C(n4_adj_85), 
         .D(n31628), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_adj_160 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [4]), 
         .Z(n29038)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_160.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_161 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [5]), 
         .Z(n29039)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_161.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_162 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [6]), 
         .Z(n29040)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_162.init = 16'h8080;
    LUT4 Select_4285_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[9]), .D(rw), .Z(n2_adj_22)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4285_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4288_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[8]), .D(rw), .Z(n2_adj_23)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4288_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_163 (.A(n1473[3]), .B(n31453), .C(\buffer[4] [7]), 
         .Z(n29041)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_163.init = 16'h8080;
    LUT4 Select_4289_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[7]), .D(rw), .Z(n3)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4289_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_164 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [0]), 
         .Z(n29042)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_164.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_165 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [1]), 
         .Z(n29043)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_165.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_166 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [2]), 
         .Z(n29044)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_166.init = 16'h8080;
    LUT4 i2_4_lut_adj_167 (.A(databus[18]), .B(n5_adj_88), .C(n1473[13]), 
         .D(n29036), .Z(n27543)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_167.init = 16'hffec;
    LUT4 select_2129_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1473[4]), 
         .C(rx_data[2]), .D(n29360), .Z(n5_adj_88)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_168 (.A(databus[19]), .B(n5_adj_89), .C(n1473[13]), 
         .D(n29037), .Z(n27533)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_168.init = 16'hffec;
    LUT4 Select_4290_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[6]), .D(rw), .Z(n3_adj_24)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4290_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4291_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[5]), .D(rw), .Z(n3_adj_25)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4291_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_169 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [3]), 
         .Z(n29045)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_169.init = 16'h8080;
    LUT4 sendcount_1__bdd_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(sendcount[3]), 
         .D(sendcount[2]), .Z(n30822)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_1__bdd_4_lut.init = 16'h6aaa;
    LUT4 select_2129_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1473[4]), 
         .C(rx_data[3]), .D(n29360), .Z(n5_adj_89)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_333_3_lut_4_lut (.A(register_addr[3]), .B(n31595), 
         .C(register_addr[2]), .D(n31589), .Z(n31476)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_333_3_lut_4_lut.init = 16'hfffe;
    LUT4 Select_4292_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[4]), .D(rw), .Z(n3_adj_26)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4292_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4293_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[3]), .D(rw), .Z(n3_adj_27)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4293_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4294_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[2]), .D(rw), .Z(n3_adj_28)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4294_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_170 (.A(databus[20]), .B(n5_adj_95), .C(n1473[13]), 
         .D(n29038), .Z(n27426)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_170.init = 16'hffec;
    LUT4 Select_4295_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[1]), .D(rw), .Z(n3_adj_29)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4295_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 select_2129_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1473[4]), 
         .C(rx_data[4]), .D(n29360), .Z(n5_adj_95)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 sendcount_4__bdd_3_lut (.A(sendcount[4]), .B(n30822), .C(\sendcount[1] ), 
         .Z(n30823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_171 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [4]), 
         .Z(n29014)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_171.init = 16'h8080;
    LUT4 i2_4_lut_adj_172 (.A(databus[21]), .B(n5_adj_97), .C(n1473[13]), 
         .D(n29039), .Z(n27478)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_172.init = 16'hffec;
    LUT4 select_2129_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1473[4]), 
         .C(rx_data[5]), .D(n29360), .Z(n5_adj_97)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_173 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [5]), 
         .Z(n29017)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_173.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_174 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [6]), 
         .Z(n29015)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_174.init = 16'h8080;
    LUT4 i2_4_lut_adj_175 (.A(databus[22]), .B(n5_adj_98), .C(n1473[13]), 
         .D(n29040), .Z(n27610)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_175.init = 16'hffec;
    LUT4 Select_4296_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[0]), .D(rw), .Z(n3_adj_30)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4296_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 select_2129_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1473[4]), 
         .C(rx_data[6]), .D(n29360), .Z(n5_adj_98)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4219_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[31]), .D(rw), .Z(n2_adj_31)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4219_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_176 (.A(n1473[3]), .B(n31453), .C(\buffer[5] [7]), 
         .Z(n29016)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_176.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_177 (.A(n1473[4]), .B(n31552), .C(bufcount[0]), 
         .D(n31450), .Z(n27625)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_177.init = 16'hd222;
    LUT4 Select_4222_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[30]), .D(rw), .Z(n2_adj_32)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4222_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_178 (.A(databus[23]), .B(n5_adj_102), .C(n1473[13]), 
         .D(n29041), .Z(n27496)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_178.init = 16'hffec;
    LUT4 select_2129_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1473[4]), 
         .C(rx_data[7]), .D(n29360), .Z(n5_adj_102)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_179 (.A(databus[24]), .B(n5_adj_103), .C(n1473[13]), 
         .D(n29042), .Z(n27513)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_179.init = 16'hffec;
    LUT4 select_2129_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1473[4]), 
         .C(rx_data[0]), .D(n29361), .Z(n5_adj_103)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4225_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[29]), .D(rw), .Z(n2_adj_33)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4225_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4228_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[28]), .D(rw), .Z(n2_adj_34)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4228_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4231_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[27]), .D(rw), .Z(n2_adj_35)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4231_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_180 (.A(databus[25]), .B(n5_adj_107), .C(n1473[13]), 
         .D(n29043), .Z(n27512)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_180.init = 16'hffec;
    LUT4 Select_4234_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31507), 
         .C(read_value[26]), .D(rw), .Z(n2_adj_36)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4234_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i17815_3_lut_4_lut (.A(n31500), .B(n31599), .C(n57_adj_109), 
         .D(escape), .Z(n10974)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i17815_3_lut_4_lut.init = 16'h7780;
    LUT4 select_2129_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1473[4]), 
         .C(rx_data[1]), .D(n29361), .Z(n5_adj_107)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_335_3_lut_4_lut (.A(n31595), .B(register_addr[5]), 
         .C(prev_select_adj_6), .D(n31544), .Z(n31478)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_335_3_lut_4_lut.init = 16'hfffb;
    LUT4 mux_1553_i12_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[11]), 
         .D(n224[11]), .Z(n3921[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_339_3_lut_4_lut (.A(n31595), .B(register_addr[5]), 
         .C(\select[4] ), .D(n31544), .Z(n31482)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_rep_339_3_lut_4_lut.init = 16'h0040;
    LUT4 mux_1553_i19_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[18]), 
         .D(n224[18]), .Z(n3921[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i18_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[17]), 
         .D(n224[17]), .Z(n3921[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_181 (.A(databus[26]), .B(n5_adj_110), .C(n1473[13]), 
         .D(n29044), .Z(n27476)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_181.init = 16'hffec;
    LUT4 i1_2_lut_rep_360_3_lut_4_lut (.A(register_addr[4]), .B(n31555), 
         .C(n31595), .D(register_addr[5]), .Z(n31503)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_360_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_364_3_lut_4_lut (.A(register_addr[4]), .B(n31555), 
         .C(register_addr[5]), .D(n31595), .Z(n31507)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_364_3_lut_4_lut.init = 16'hffef;
    LUT4 select_2129_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1473[4]), 
         .C(rx_data[2]), .D(n29361), .Z(n5_adj_110)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 i24_3_lut_4_lut_adj_182 (.A(bufcount[0]), .B(n31553), .C(\buffer[1] [0]), 
         .D(rx_data[0]), .Z(n11_adj_111)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_182.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_183 (.A(bufcount[0]), .B(n31553), .C(rx_data[1]), 
         .D(\buffer[1] [1]), .Z(n11_adj_112)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_183.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_184 (.A(bufcount[0]), .B(n31553), .C(rx_data[2]), 
         .D(\buffer[1] [2]), .Z(n11_adj_113)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_184.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_185 (.A(bufcount[0]), .B(n31553), .C(\buffer[1] [3]), 
         .D(rx_data[3]), .Z(n11_adj_114)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_185.init = 16'hf2d0;
    LUT4 i2_4_lut_adj_186 (.A(databus[27]), .B(n5_adj_115), .C(n1473[13]), 
         .D(n29045), .Z(n27511)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_186.init = 16'hffec;
    LUT4 i2_3_lut_4_lut_adj_187 (.A(register_addr[1]), .B(n31476), .C(register_addr[0]), 
         .D(n14453), .Z(n9537)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_187.init = 16'h2000;
    LUT4 n31453_bdd_4_lut_23119 (.A(n31453), .B(n31551), .C(n1473[0]), 
         .D(n1473[3]), .Z(n31949)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n31453_bdd_4_lut_23119.init = 16'hee0f;
    LUT4 i24_3_lut_4_lut_adj_188 (.A(bufcount[0]), .B(n31553), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_116)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_188.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_189 (.A(bufcount[0]), .B(n31553), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_117)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_189.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_190 (.A(bufcount[0]), .B(n31553), .C(rx_data[6]), 
         .D(\buffer[1] [6]), .Z(n11_adj_118)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_190.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_191 (.A(bufcount[0]), .B(n31553), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_119)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_191.init = 16'hf2d0;
    LUT4 select_2129_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1473[4]), 
         .C(rx_data[3]), .D(n29361), .Z(n5_adj_115)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_279 (.A(register_addr[4]), .B(n35), .Z(n31422)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_279.init = 16'h8888;
    LUT4 mux_1553_i17_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[16]), 
         .D(n224[16]), .Z(n3921[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_192 (.A(databus[28]), .B(n5_adj_120), .C(n1473[13]), 
         .D(n29014), .Z(n27510)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_192.init = 16'hffec;
    FD1P3IX send_491 (.D(n33383), .SP(n2224), .CD(n27464), .CK(debug_c_c), 
            .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 select_2129_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1473[4]), 
         .C(rx_data[4]), .D(n29361), .Z(n5_adj_120)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_193 (.A(databus[29]), .B(n5_adj_121), .C(n1473[13]), 
         .D(n29017), .Z(n27465)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_193.init = 16'hffec;
    LUT4 i4_2_lut_rep_405 (.A(n1491), .B(n1473[15]), .Z(n31548)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_405.init = 16'heeee;
    LUT4 select_2129_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1473[4]), 
         .C(rx_data[5]), .D(n29361), .Z(n5_adj_121)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_369_3_lut (.A(n1491), .B(n1473[15]), .C(n1473[12]), 
         .Z(n31512)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_369_3_lut.init = 16'hfefe;
    LUT4 i507_2_lut (.A(n1473[3]), .B(n1473[4]), .Z(n1874)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i507_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_rep_406 (.A(n1473[19]), .B(n1473[3]), .C(n1473[11]), 
         .Z(n31549)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_rep_406.init = 16'hfefe;
    LUT4 i3_2_lut_4_lut (.A(n1473[19]), .B(n1473[3]), .C(n1473[11]), .D(n31550), 
         .Z(n9_adj_122)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_194 (.A(databus[30]), .B(n5_adj_123), .C(n1473[13]), 
         .D(n29015), .Z(n27505)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_194.init = 16'hffec;
    LUT4 select_2129_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1473[4]), 
         .C(rx_data[6]), .D(n29361), .Z(n5_adj_123)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i2_3_lut_rep_407 (.A(n1473[7]), .B(n1473[13]), .C(n1473[5]), 
         .Z(n31550)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_407.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(n1473[7]), .B(n1473[13]), .C(n1473[5]), .D(n1473[6]), 
         .Z(n6)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1553_i11_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[10]), 
         .D(n224[10]), .Z(n3921[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_195 (.A(databus[31]), .B(n5_adj_124), .C(n1473[13]), 
         .D(n29016), .Z(n27499)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_195.init = 16'hffec;
    LUT4 select_2129_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1473[4]), 
         .C(rx_data[7]), .D(n29361), .Z(n5_adj_124)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 n31453_bdd_4_lut (.A(bufcount[1]), .B(n1473[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n31951)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n31453_bdd_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_302_3_lut_4_lut (.A(n31555), .B(n31514), .C(\select[4] ), 
         .D(register_addr[5]), .Z(n31445)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_302_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_408 (.A(debug_c_7), .B(escape), .Z(n31551)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_408.init = 16'hdddd;
    LUT4 i2_3_lut_rep_307_4_lut (.A(debug_c_7), .B(escape), .C(n31453), 
         .D(n1473[4]), .Z(n31450)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i2_3_lut_rep_307_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_196 (.A(n31555), .B(n31514), .C(\read_size[2] ), 
         .D(register_addr[5]), .Z(n29234)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_196.init = 16'h0040;
    LUT4 i1_2_lut_rep_301_3_lut_4_lut (.A(n31555), .B(n31514), .C(register_addr[5]), 
         .D(\select[4] ), .Z(n31444)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_301_3_lut_4_lut.init = 16'h4000;
    LUT4 i15596_3_lut_rep_409 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n31552)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15596_3_lut_rep_409.init = 16'hecec;
    LUT4 i2_2_lut_rep_398_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1473[4]), .Z(n31541)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_398_4_lut.init = 16'hecff;
    LUT4 i1_2_lut_4_lut_adj_197 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1473[4]), .Z(n7_adj_125)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_197.init = 16'hec00;
    LUT4 equal_201_i4_2_lut_rep_410 (.A(bufcount[1]), .B(bufcount[2]), .Z(n31553)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam equal_201_i4_2_lut_rep_410.init = 16'heeee;
    LUT4 mux_1553_i16_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[15]), 
         .D(n224[15]), .Z(n3921[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i15_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[14]), 
         .D(n224[14]), .Z(n3921[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i2937_2_lut_rep_379_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n31522)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i2937_2_lut_rep_379_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_198 (.A(n31544), .B(n31532), .C(n33384), 
         .D(\select[4] ), .Z(n52)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_198.init = 16'h1000;
    LUT4 i1_4_lut_adj_199 (.A(n1473[4]), .B(\buffer[0] [1]), .C(n11_adj_44), 
         .D(n14_c), .Z(n28666)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_199.init = 16'heca0;
    LUT4 i1_4_lut_adj_200 (.A(n1473[4]), .B(\buffer[0] [2]), .C(n11_adj_45), 
         .D(n14_c), .Z(n28658)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_200.init = 16'heca0;
    LUT4 i1_2_lut_rep_299_3_lut_4_lut (.A(n31544), .B(n31532), .C(prev_select_adj_5), 
         .D(\select[4] ), .Z(n31442)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_299_3_lut_4_lut.init = 16'h0100;
    LUT4 mux_1553_i14_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[13]), 
         .D(n224[13]), .Z(n3921[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i15591_1_lut_3_lut_4_lut (.A(n31589), .B(n31538), .C(n29236), 
         .D(register_addr[2]), .Z(n176)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i15591_1_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i1_2_lut_3_lut_4_lut_adj_201 (.A(rw), .B(n31448), .C(register_addr[0]), 
         .D(n31570), .Z(n16012)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_201.init = 16'h1000;
    LUT4 i15590_3_lut_rep_313_4_lut (.A(n31589), .B(n31538), .C(n29236), 
         .D(register_addr[2]), .Z(n31456)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i15590_3_lut_rep_313_4_lut.init = 16'hfeee;
    LUT4 i22017_2_lut (.A(esc_data[5]), .B(esc_data[6]), .Z(n29573)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22017_2_lut.init = 16'heeee;
    LUT4 i22360_2_lut_3_lut_4_lut (.A(rw), .B(n31448), .C(register_addr[0]), 
         .D(n31581), .Z(n13907)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i22360_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i21901_2_lut_rep_412 (.A(register_addr[2]), .B(register_addr[3]), 
         .Z(n31555)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21901_2_lut_rep_412.init = 16'heeee;
    LUT4 i4460_2_lut_3_lut_4_lut (.A(rw), .B(n31448), .C(register_addr[0]), 
         .D(n31581), .Z(n11235)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4460_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_291_3_lut_4_lut (.A(n31589), .B(n31538), .C(register_addr[1]), 
         .D(register_addr[2]), .Z(n31434)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_291_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_202 (.A(n1473[4]), .B(\buffer[0] [3]), .C(n11_adj_46), 
         .D(n14_c), .Z(n28616)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_202.init = 16'heca0;
    LUT4 n30304_bdd_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n30304), .D(n31523), .Z(n30305)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n30304_bdd_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_1553_i10_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[9]), 
         .D(n224[9]), .Z(n3921[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 esc_data_1__bdd_4_lut (.A(esc_data[1]), .B(esc_data[3]), .C(esc_data[2]), 
         .D(esc_data[4]), .Z(n30339)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)))+!A (B+(C+(D)))) */ ;
    defparam esc_data_1__bdd_4_lut.init = 16'hd7fe;
    LUT4 i1_2_lut_adj_203 (.A(rx_data[4]), .B(rx_data[1]), .Z(n29276)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_203.init = 16'h8888;
    LUT4 mux_1553_i1_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[0]), 
         .D(n224[0]), .Z(n3921[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i32_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[31]), 
         .D(n224[31]), .Z(n3921[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_4_lut_adj_204 (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n28), .D(n31523), .Z(n29220)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_3_lut_4_lut_adj_204.init = 16'h0010;
    LUT4 mux_1553_i31_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[30]), 
         .D(n224[30]), .Z(n3921[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_305_3_lut_4_lut (.A(n31589), .B(n31538), .C(register_addr[1]), 
         .D(register_addr[2]), .Z(n31448)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_305_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21962_2_lut_rep_382_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .Z(n31525)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i21962_2_lut_rep_382_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_276_3_lut_4_lut (.A(register_addr[4]), .B(n31540), 
         .C(n29230), .D(n31595), .Z(n31419)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_276_3_lut_4_lut.init = 16'h0010;
    LUT4 n30302_bdd_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n30302), .D(n31523), .Z(n30303)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n30302_bdd_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_205 (.A(register_addr[0]), .B(\control_reg[7] ), .Z(n1)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_205.init = 16'h4444;
    LUT4 i1_4_lut_adj_206 (.A(n1473[4]), .B(\buffer[0] [4]), .C(n11_adj_47), 
         .D(n14_c), .Z(n28614)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_206.init = 16'heca0;
    LUT4 i2_3_lut_rep_386_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n31595), .D(n29169), .Z(n31529)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_386_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_207 (.A(n1473[4]), .B(\buffer[0] [5]), .C(n11_adj_48), 
         .D(n14_c), .Z(n28618)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_207.init = 16'heca0;
    LUT4 i1_4_lut_adj_208 (.A(n1473[4]), .B(\buffer[0] [6]), .C(n11_adj_49), 
         .D(n14_c), .Z(n28620)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_208.init = 16'heca0;
    LUT4 i1_4_lut_adj_209 (.A(n1473[4]), .B(\buffer[0] [7]), .C(n11_adj_50), 
         .D(n14_c), .Z(n28662)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_209.init = 16'heca0;
    LUT4 i1_2_lut_rep_396_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[4]), .Z(n31539)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_396_3_lut.init = 16'h1010;
    PFUMX i8907 (.BLUT(n15678), .ALUT(n1869[1]), .C0(n1874), .Z(n15679));
    LUT4 i1_4_lut_adj_210 (.A(sendcount[4]), .B(n1_adj_126), .C(n6_adj_127), 
         .D(n13155), .Z(n9_adj_53)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_210.init = 16'hfeff;
    LUT4 equal_63_i1_4_lut (.A(sendcount[0]), .B(n13), .C(n18), .D(n14), 
         .Z(n1_adj_126)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_63_i1_4_lut.init = 16'h5556;
    LUT4 i1_4_lut_adj_211 (.A(n1473[4]), .B(\buffer[1] [0]), .C(n11_adj_111), 
         .D(n14_c), .Z(n28612)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_211.init = 16'heca0;
    LUT4 i14916_2_lut (.A(bufcount[1]), .B(n1473[0]), .Z(n15678)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14916_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_212 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n31587), .Z(n6_adj_127)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_212.init = 16'he7de;
    LUT4 i1_2_lut_3_lut_4_lut_adj_213 (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n31595), .D(register_addr[4]), .Z(n31496)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_213.init = 16'h0100;
    LUT4 i1_4_lut_adj_214 (.A(n1473[4]), .B(\buffer[1] [1]), .C(n11_adj_112), 
         .D(n14_c), .Z(n28660)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_214.init = 16'heca0;
    PFUMX i9010 (.BLUT(n15781), .ALUT(n27625), .C0(n1874), .Z(n15782));
    LUT4 i1_2_lut_rep_363_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[4]), .D(n31590), .Z(n31506)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_363_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_215 (.A(n1473[4]), .B(\buffer[1] [2]), .C(n11_adj_113), 
         .D(n14_c), .Z(n28624)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_215.init = 16'heca0;
    LUT4 i1_2_lut_rep_401_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[4]), .Z(n31544)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_401_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_216 (.A(n1473[4]), .B(\buffer[1] [3]), .C(n11_adj_114), 
         .D(n14_c), .Z(n28608)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_216.init = 16'heca0;
    LUT4 i1_4_lut_adj_217 (.A(n1473[4]), .B(\buffer[1] [4]), .C(n11_adj_116), 
         .D(n14_c), .Z(n28610)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_217.init = 16'heca0;
    LUT4 n29161_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n30340)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n29161_bdd_4_lut.init = 16'h4001;
    LUT4 mux_1553_i30_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[29]), 
         .D(n224[29]), .Z(n3921[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_218 (.A(n1473[4]), .B(\buffer[1] [5]), .C(n11_adj_117), 
         .D(n14_c), .Z(n28586)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_218.init = 16'heca0;
    LUT4 i1_4_lut_adj_219 (.A(n1473[4]), .B(\buffer[1] [6]), .C(n11_adj_118), 
         .D(n14_c), .Z(n28622)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_219.init = 16'heca0;
    LUT4 mux_1553_i29_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[28]), 
         .D(n224[28]), .Z(n3921[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_220 (.A(n1473[4]), .B(\buffer[1] [7]), .C(n11_adj_119), 
         .D(n14_c), .Z(n28606)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_220.init = 16'heca0;
    LUT4 i2_4_lut_adj_221 (.A(databus[0]), .B(n5_adj_130), .C(n1473[13]), 
         .D(n29018), .Z(n27601)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_221.init = 16'hffec;
    LUT4 select_2129_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1473[4]), 
         .C(rx_data[0]), .D(n29357), .Z(n5_adj_130)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_222 (.A(databus[1]), .B(n5_adj_131), .C(n1473[13]), 
         .D(n29019), .Z(n27599)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_222.init = 16'hffec;
    LUT4 mux_1553_i9_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[8]), 
         .D(n224[8]), .Z(n3921[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i28_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[27]), 
         .D(n224[27]), .Z(n3921[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 select_2129_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1473[4]), 
         .C(rx_data[1]), .D(n29357), .Z(n5_adj_131)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2129_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i14921_2_lut_3_lut (.A(n1473[0]), .B(n1473[8]), .C(\select[7] ), 
         .Z(n15666)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14921_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_3_lut (.A(n27441), .B(\control_reg[7]_adj_37 ), .C(n31600), 
         .Z(n32)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut.init = 16'h0808;
    LUT4 mux_1553_i8_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[7]), 
         .D(n224[7]), .Z(n3921[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i14919_2_lut_3_lut (.A(n1473[0]), .B(n1473[8]), .C(\select[5] ), 
         .Z(n15670)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14919_2_lut_3_lut.init = 16'h1010;
    LUT4 i957_2_lut (.A(n1473[5]), .B(n31500), .Z(n2807)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i957_2_lut.init = 16'h8888;
    LUT4 i15119_2_lut_3_lut (.A(n1473[0]), .B(n1473[8]), .C(\select[2] ), 
         .Z(n16684)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15119_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_223 (.A(n1473[0]), .B(n1473[8]), .C(\select[4] ), 
         .Z(n15674)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_223.init = 16'h1010;
    LUT4 i1_2_lut_adj_224 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_224.init = 16'h4444;
    LUT4 i2_4_lut_adj_225 (.A(databus[2]), .B(n5), .C(n1473[13]), .D(n29020), 
         .Z(n27602)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_225.init = 16'hffec;
    LUT4 mux_1895_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n5833), 
         .Z(n5824[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1895_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_85)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_rep_427 (.A(\select[5] ), .B(prev_select_adj_38), .Z(n31570)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_427.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\select[5] ), .B(prev_select_adj_38), 
         .C(\reset_count[14] ), .D(n22483), .Z(n2869)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_1553_i7_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[6]), 
         .D(n224[6]), .Z(n3921[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i6_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[5]), 
         .D(n224[5]), .Z(n3921[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i8_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[7]), 
         .D(n224_adj_91[7]), .Z(n4094[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i7_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[6]), 
         .D(n224_adj_91[6]), .Z(n4094[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i14929_2_lut (.A(bufcount[0]), .B(n1473[0]), .Z(n15781)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14929_2_lut.init = 16'h2222;
    LUT4 mux_1553_i5_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[4]), 
         .D(n224[4]), .Z(n3921[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i4_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[3]), 
         .D(n224[3]), .Z(n3921[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_432 (.A(rw), .B(register_addr[5]), .Z(n31575)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_432.init = 16'h4444;
    LUT4 i1_2_lut_rep_271_3_lut_4_lut_4_lut (.A(n33384), .B(register_addr[5]), 
         .C(prev_select), .D(n31465), .Z(n31414)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_271_3_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 Select_4289_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31465), 
         .C(\read_value[7]_adj_71 ), .D(n33384), .Z(n2_adj_72)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4289_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1895_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n5833), 
         .Z(n5824[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1895_i3_3_lut.init = 16'hcaca;
    LUT4 Select_4291_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31465), 
         .C(\read_value[5]_adj_73 ), .D(rw), .Z(n2_adj_74)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4291_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1S3JX state_FSM_i1 (.D(n13788), .CK(debug_c_c), .PD(n31472), .Q(n1473[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_64)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i955_3_lut (.A(n1473[5]), .B(n31500), .C(n1473[10]), .Z(n2805)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i955_3_lut.init = 16'hc8c8;
    LUT4 mux_1895_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n5833), 
         .Z(n5824[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1895_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_437 (.A(n1491), .B(sendcount[4]), .Z(n31580)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_437.init = 16'h2222;
    LUT4 motor_pwm_r_c_15_bdd_2_lut_22585_3_lut (.A(n1491), .B(sendcount[4]), 
         .C(n30340), .Z(n30341)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam motor_pwm_r_c_15_bdd_2_lut_22585_3_lut.init = 16'h2020;
    LUT4 Select_4292_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31465), 
         .C(\read_value[4]_adj_75 ), .D(rw), .Z(n2_adj_76)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4292_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_adj_63)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    PFUMX i9913 (.BLUT(n16684), .ALUT(n27433), .C0(n1926), .Z(n16685));
    PFUMX i8895 (.BLUT(n15666), .ALUT(n27681), .C0(n1926), .Z(n15667));
    LUT4 mux_1598_i20_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[19]), 
         .D(n224_adj_91[19]), .Z(n4094[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_521_i5_3_lut (.A(n2746), .B(esc_data[4]), .C(n1473[18]), 
         .Z(n2215[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_521_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_226 (.A(n1473[15]), .B(n7), .C(n30733), .D(n29573), 
         .Z(n2746)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_226.init = 16'h0020;
    LUT4 Select_4290_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31465), 
         .C(\read_value[6]_adj_77 ), .D(n33384), .Z(n2_adj_78)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4290_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1553_i3_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[2]), 
         .D(n224[2]), .Z(n3921[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_440 (.A(sendcount[0]), .B(\sendcount[1] ), .Z(n31583)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_2_lut_rep_440.init = 16'h8888;
    LUT4 Select_4293_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31465), 
         .C(\read_value[3]_adj_79 ), .D(rw), .Z(n2_adj_80)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4293_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1553_i2_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[1]), 
         .D(n224[1]), .Z(n3921[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i14820_3_lut_4_lut (.A(sendcount[0]), .B(\sendcount[1] ), .C(n9_adj_53), 
         .D(sendcount[2]), .Z(n17[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i14820_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i14748_2_lut_rep_441 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n31584)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14748_2_lut_rep_441.init = 16'heeee;
    LUT4 i2_2_lut (.A(esc_data[7]), .B(esc_data[0]), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_391_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n31534)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_391_3_lut.init = 16'h1e1e;
    LUT4 i3395_2_lut_rep_442 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n31585)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i3395_2_lut_rep_442.init = 16'h9999;
    LUT4 Select_4294_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31465), 
         .C(\read_value[2]_adj_81 ), .D(rw), .Z(n2_adj_82)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4294_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4296_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31465), 
         .C(\read_value[0]_adj_83 ), .D(n33384), .Z(n2_adj_84)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4296_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_521_i4_3_lut (.A(n2746), .B(esc_data[3]), .C(n1473[18]), 
         .Z(n2215[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_521_i4_3_lut.init = 16'hcaca;
    PFUMX i22641 (.BLUT(n30706), .ALUT(n13_adj_151), .C0(n5833), .Z(n30707));
    LUT4 mux_521_i2_3_lut (.A(n2746), .B(esc_data[1]), .C(n1473[18]), 
         .Z(n2215[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_521_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1598_i1_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[0]), 
         .D(n224_adj_91[0]), .Z(n4094[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i19_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[18]), 
         .D(n224_adj_91[18]), .Z(n4094[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i14821_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_adj_53), .Z(n17[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i14821_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 n13157_bdd_4_lut_22663_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n30705)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n13157_bdd_4_lut_22663_4_lut.init = 16'h6420;
    LUT4 mux_1598_i32_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[31]), 
         .D(n224_adj_91[31]), .Z(n4094[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_521_i1_3_lut (.A(n2746), .B(esc_data[0]), .C(n1473[18]), 
         .Z(n2215[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_521_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_adj_227 (.A(n27444), .B(\control_reg[7] ), .C(n31600), 
         .Z(n34)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_227.init = 16'h0808;
    LUT4 i3_4_lut (.A(register_addr[1]), .B(register_addr[2]), .C(n31538), 
         .D(n29255), .Z(n29256)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_4_lut.init = 16'h0200;
    LUT4 mux_1553_i21_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[20]), 
         .D(n224[20]), .Z(n3921[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i18_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[17]), 
         .D(n224_adj_91[17]), .Z(n4094[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i31_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[30]), 
         .D(n224_adj_91[30]), .Z(n4094[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i27_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[26]), 
         .D(n224[26]), .Z(n3921[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i4437_3_lut (.A(n1473[19]), .B(n1473[18]), .C(busy), .Z(n11202)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4437_3_lut.init = 16'hcece;
    LUT4 i3_3_lut_4_lut (.A(n31427), .B(n31575), .C(n31496), .D(n19331), 
         .Z(n9330)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_1553_i26_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[25]), 
         .D(n224[25]), .Z(n3921[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i26_3_lut_4_lut.init = 16'hf780;
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2805), .CK(debug_c_c), 
            .Q(register_addr[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 i5581_3_lut (.A(busy), .B(n1485), .C(n1473[19]), .Z(n12349)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5581_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut_adj_228 (.A(sendcount[0]), .B(sendcount[3]), .Z(n13_adj_151)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_228.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_446 (.A(register_addr[5]), .B(register_addr[4]), .Z(n31589)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_446.init = 16'heeee;
    LUT4 i12432_3_lut (.A(\register[0][5] ), .B(expansion5_c), .C(register_addr[1]), 
         .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i12432_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_229 (.A(register_addr[1]), .B(\register[1][5] ), .Z(n159)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_229.init = 16'h4444;
    LUT4 i1_2_lut_adj_230 (.A(n1473[6]), .B(n1473[11]), .Z(n1926)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_230.init = 16'heeee;
    LUT4 i5_4_lut (.A(n9_adj_122), .B(n1473[15]), .C(n8), .D(n1473[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_adj_231 (.A(n1488), .B(n1473[9]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut_adj_231.init = 16'heeee;
    LUT4 i1_4_lut_adj_232 (.A(n31548), .B(n1473[7]), .C(n10_adj_157), 
         .D(n31549), .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_232.init = 16'hfffe;
    LUT4 reduce_or_2658_i1_2_lut_3_lut_4_lut_4_lut (.A(n31477), .B(register_addr[0]), 
         .C(n31476), .D(register_addr[1]), .Z(n9378)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;
    defparam reduce_or_2658_i1_2_lut_3_lut_4_lut_4_lut.init = 16'h555d;
    LUT4 i1_2_lut_rep_362_3_lut_4_lut (.A(register_addr[5]), .B(register_addr[4]), 
         .C(n31595), .D(register_addr[3]), .Z(n31505)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_362_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4_4_lut (.A(n1473[2]), .B(n1473[10]), .C(n1473[18]), .D(n1473[6]), 
         .Z(n10_adj_157)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_233 (.A(\buffer[0] [3]), .B(\buffer[0] [5]), .C(\buffer[0] [4]), 
         .D(\buffer[0] [6]), .Z(n28916)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i3_4_lut_adj_233.init = 16'hfffe;
    LUT4 i1_2_lut_rep_272_3_lut_4_lut (.A(\select[4] ), .B(n31469), .C(n29491), 
         .D(prev_select_adj_85), .Z(n31415)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_272_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_adj_234 (.A(register_addr[1]), .B(\steps_reg[7] ), .Z(n11)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_234.init = 16'h8888;
    LUT4 i4_4_lut_adj_235 (.A(n1473[4]), .B(n31512), .C(n1485), .D(n6), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_235.init = 16'hfffe;
    LUT4 mux_1598_i17_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[16]), 
         .D(n224_adj_91[16]), .Z(n4094[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i6_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[5]), 
         .D(n224_adj_91[5]), .Z(n4094[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i16_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[15]), 
         .D(n224_adj_91[15]), .Z(n4094[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i22013_2_lut_rep_452 (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .Z(n31595)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22013_2_lut_rep_452.init = 16'heeee;
    LUT4 i21907_2_lut_rep_400_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[5]), .Z(n31543)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i21907_2_lut_rep_400_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_371_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[4]), .Z(n31514)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_371_3_lut.init = 16'h1010;
    LUT4 i22074_3_lut_rep_380_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[4]), .D(register_addr[5]), .Z(n31523)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22074_3_lut_rep_380_4_lut.init = 16'hfffe;
    FD1P3IX buffer_0___i2 (.D(n28666), .SP(n13041), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n28658), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n28616), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n28614), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n28618), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n28620), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n28662), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n28612), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n28660), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n28624), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n28608), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n28610), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n28586), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n28622), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n28606), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n27601), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n27599), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n27602), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n27597), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n27538), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i22 (.D(n27548), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    FD1P3IX buffer_0___i23 (.D(n27556), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n27524), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n27504), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n27472), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n27532), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n27557), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n27491), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n27555), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n27554), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n27551), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n27550), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n27500), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n27543), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n27533), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n27426), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n27478), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n27610), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n27496), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n27513), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n27512), .SP(n9471), .CD(n31472), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n27476), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n27511), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n27510), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n27465), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n27505), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n27499), .SP(n9471), .CD(n33389), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_389_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[5]), .Z(n31532)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_389_3_lut.init = 16'hfefe;
    LUT4 i4384_2_lut_rep_358_3_lut_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[4]), .D(register_addr[5]), .Z(n31501)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i4384_2_lut_rep_358_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_395_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[3]), .Z(n31538)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_395_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_236 (.A(n45_adj_163), .B(n112), .C(register_addr[0]), 
         .D(n28899), .Z(n6005)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_236.init = 16'h333b;
    LUT4 i1_2_lut_3_lut_adj_237 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29360)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_237.init = 16'hfbfb;
    LUT4 i18000_3_lut (.A(n31600), .B(\register[2] [0]), .C(register_addr[1]), 
         .Z(n45_adj_163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i18000_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_238 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29361)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_238.init = 16'hbfbf;
    LUT4 i4_4_lut_adj_239 (.A(n1473[11]), .B(n1473[8]), .C(n1473[13]), 
         .D(n1473[10]), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_239.init = 16'hfffe;
    LUT4 i1_2_lut_adj_240 (.A(register_addr[1]), .B(\steps_reg[5] ), .Z(n14_adj_86)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_240.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_241 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29357)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_241.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_242 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29358)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_242.init = 16'hbfbf;
    LUT4 mux_1598_i15_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[14]), 
         .D(n224_adj_91[14]), .Z(n4094[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i14_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[13]), 
         .D(n224_adj_91[13]), .Z(n4094[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i37_3_lut (.A(\register[0][4] ), .B(expansion4_out), .C(register_addr[1]), 
         .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i37_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_456 (.A(n1473[3]), .B(debug_c_7), .Z(n31599)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_456.init = 16'h8888;
    LUT4 i1_2_lut_adj_243 (.A(register_addr[1]), .B(\register[1][4] ), .Z(n19)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_adj_243.init = 16'h4444;
    LUT4 mux_1598_i5_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[4]), 
         .D(n224_adj_91[4]), .Z(n4094[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_rep_457 (.A(force_pause), .B(\register[0][2] ), .C(timeout_pause), 
         .Z(n31600)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[6:17])
    defparam i2_3_lut_rep_457.init = 16'hfefe;
    LUT4 mux_1598_i4_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[3]), 
         .D(n224_adj_91[3]), .Z(n4094[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i3_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[2]), 
         .D(n224_adj_91[2]), .Z(n4094[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_244 (.A(register_addr[1]), .B(\steps_reg[6] ), .Z(n13_adj_87)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_244.init = 16'h8888;
    LUT4 i15237_2_lut_rep_393_4_lut (.A(force_pause), .B(\register[0][2] ), 
         .C(timeout_pause), .D(\register[0][7] ), .Z(n31536)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[6:17])
    defparam i15237_2_lut_rep_393_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_4_lut_adj_245 (.A(force_pause), .B(\register[0][2] ), 
         .C(timeout_pause), .D(clk_1Hz), .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[6:17])
    defparam i1_2_lut_4_lut_adj_245.init = 16'hfffe;
    LUT4 i22318_2_lut_2_lut (.A(n31500), .B(n13041), .Z(n9471)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22318_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_1598_i2_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[1]), 
         .D(n224_adj_91[1]), .Z(n4094[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_246 (.A(register_addr[1]), .B(\steps_reg[3] ), .Z(n12)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_246.init = 16'h8888;
    LUT4 i22_3_lut (.A(\control_reg[4] ), .B(\div_factor_reg[4] ), .C(register_addr[1]), 
         .Z(n12_adj_172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i22_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_247 (.A(register_addr[1]), .B(\steps_reg[4] ), .Z(n6_adj_173)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_adj_247.init = 16'h8888;
    LUT4 i1_4_lut_adj_248 (.A(n29162), .B(debug_c_7), .C(n1473[0]), .D(n1473[1]), 
         .Z(n13788)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_248.init = 16'hbbba;
    LUT4 i3_4_lut_adj_249 (.A(sendcount[3]), .B(n31584), .C(sendcount[2]), 
         .D(n31580), .Z(n29162)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_249.init = 16'h0200;
    LUT4 i1_2_lut_adj_250 (.A(register_addr[0]), .B(\control_reg[7]_adj_88 ), 
         .Z(n8635)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_250.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_251 (.A(n31570), .B(n31423), .C(register_addr[0]), 
         .D(n31511), .Z(n13947)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_251.init = 16'h0f02;
    LUT4 i1_2_lut_3_lut_4_lut_adj_252 (.A(n31570), .B(n31423), .C(register_addr[0]), 
         .D(n31511), .Z(n12368)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_252.init = 16'hf020;
    LUT4 mux_1598_i13_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[12]), 
         .D(n224_adj_91[12]), .Z(n4094[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i23_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[22]), 
         .D(n224[22]), .Z(n3921[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 i21939_2_lut (.A(n33384), .B(register_addr[5]), .Z(n29491)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21939_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_253 (.A(prev_select_adj_85), .B(n29169), .C(n29491), 
         .D(n31465), .Z(n9300)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut_adj_253.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_254 (.A(n31595), .B(n31506), .C(n31511), 
         .D(n29230), .Z(n14522)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_254.init = 16'hf1f0;
    FD1S3IX state_FSM_i2 (.D(n28692), .CK(debug_c_c), .CD(n33389), .Q(n1473[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    LUT4 i2_3_lut_adj_255 (.A(n29230), .B(n35), .C(register_addr[4]), 
         .Z(n4006)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut_adj_255.init = 16'h0808;
    LUT4 n79_bdd_4_lut (.A(n79), .B(n159), .C(register_addr[0]), .D(n31486), 
         .Z(n31406)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n79_bdd_4_lut.init = 16'h00ca;
    LUT4 i2_4_lut_adj_256 (.A(n31478), .B(register_addr[5]), .C(\select[4] ), 
         .D(rw), .Z(n29230)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_4_lut_adj_256.init = 16'h0040;
    LUT4 mux_1598_i30_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[29]), 
         .D(n224_adj_91[29]), .Z(n4094[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i30_3_lut_4_lut.init = 16'hf780;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n31468), .CD(n16769), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n31468), .CD(n16769), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n31468), .CD(n16769), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n31468), .CD(n16769), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n13833), .CD(n16767), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n13833), .CD(n16767), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n13833), .CD(n16767), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n13833), .CD(n16767), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 i2_2_lut_4_lut_4_lut (.A(n31477), .B(n31476), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n27679)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D))))) */ ;
    defparam i2_2_lut_4_lut_4_lut.init = 16'h5775;
    LUT4 i2_3_lut_adj_257 (.A(n27483), .B(\control_reg[7]_adj_88 ), .C(n31600), 
         .Z(n32_adj_89)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_257.init = 16'h0808;
    LUT4 i9992_2_lut_3_lut_4_lut_4_lut (.A(n31477), .B(n14453), .C(n31476), 
         .D(register_addr[1]), .Z(n16764)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B))) */ ;
    defparam i9992_2_lut_3_lut_4_lut_4_lut.init = 16'h4c44;
    FD1S3IX state_FSM_i3 (.D(n13464), .CK(debug_c_c), .CD(n33389), .Q(n1473[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n12481), .CK(debug_c_c), .CD(n33389), .Q(n1473[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n29228), .CK(debug_c_c), .CD(n33389), .Q(n1473[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n29204), .CK(debug_c_c), .CD(n33389), .Q(n1473[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1473[5]), .CK(debug_c_c), .CD(n33389), .Q(n1473[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1473[6]), .CK(debug_c_c), .CD(n33389), .Q(n1473[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1473[7]), .CK(debug_c_c), .CD(n33389), .Q(n1473[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1473[8]), .CK(debug_c_c), .CD(n33389), 
            .Q(n1473[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1578), .CK(debug_c_c), .CD(n33389), .Q(n1473[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1473[10]), .CK(debug_c_c), .CD(n33389), 
            .Q(n1473[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1473[11]), .CK(debug_c_c), .CD(n33389), 
            .Q(n1473[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1473[12]), .CK(debug_c_c), .CD(n33389), 
            .Q(n1473[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1584), .CK(debug_c_c), .CD(n33389), .Q(n1491));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1585), .CK(debug_c_c), .CD(n33389), .Q(n1473[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n11216), .CK(debug_c_c), .CD(n33389), .Q(n1473[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n12347), .CK(debug_c_c), .CD(n33389), .Q(n1488));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n28604), .CK(debug_c_c), .CD(n33389), .Q(n1473[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n11202), .CK(debug_c_c), .CD(n33389), .Q(n1473[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i21 (.D(n12349), .CK(debug_c_c), .CD(n33389), .Q(n1485));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    LUT4 mux_1598_i29_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[28]), 
         .D(n224_adj_91[28]), .Z(n4094[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i28_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[27]), 
         .D(n224_adj_91[27]), .Z(n4094[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i28_3_lut_4_lut.init = 16'hf780;
    FD1P3AX rw_498_rep_466 (.D(n1473[10]), .SP(n2805), .CK(debug_c_c), 
            .Q(n33384));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_466.GSR = "ENABLED";
    LUT4 mux_1598_i27_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[26]), 
         .D(n224_adj_91[26]), .Z(n4094[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i5_4_lut_adj_258 (.A(n9), .B(\select[4] ), .C(n8_adj_182), .D(register_addr[4]), 
         .Z(n9304)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i5_4_lut_adj_258.init = 16'h0080;
    LUT4 mux_1598_i26_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[25]), 
         .D(n224_adj_91[25]), .Z(n4094[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_2_lut_adj_259 (.A(register_addr[5]), .B(prev_select_adj_6), 
         .Z(n8_adj_182)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_2_lut_adj_259.init = 16'h2222;
    LUT4 i15042_3_lut_4_lut (.A(n31475), .B(n1491), .C(n9_adj_53), .D(sendcount[0]), 
         .Z(n15[0])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i15042_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i1_2_lut_adj_260 (.A(register_addr[5]), .B(register_addr[4]), .Z(n29255)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_260.init = 16'h8888;
    LUT4 i2_3_lut_rep_283_4_lut (.A(register_addr[1]), .B(n31476), .C(n31464), 
         .D(prev_select_adj_90), .Z(n31426)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_283_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut_adj_261 (.A(register_addr[0]), .B(register_addr[1]), .Z(n19331)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_261.init = 16'hbbbb;
    LUT4 mux_1598_i25_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[24]), 
         .D(n224_adj_91[24]), .Z(n4094[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_262 (.A(n31522), .B(debug_c_7), .C(n13489), .D(n8_adj_185), 
         .Z(n28692)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_262.init = 16'hdc50;
    LUT4 i1_3_lut (.A(n31453), .B(n1473[1]), .C(n1473[0]), .Z(n8_adj_185)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i4_4_lut_adj_263 (.A(n7_adj_186), .B(n29276), .C(rx_data[2]), 
         .D(rx_data[0]), .Z(n13489)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i4_4_lut_adj_263.init = 16'h8000;
    LUT4 i9991_2_lut_3_lut_4_lut_4_lut (.A(n31477), .B(n14453), .C(n31476), 
         .D(register_addr[1]), .Z(n16763)) /* synthesis lut_function=(A (B (C+!(D)))) */ ;
    defparam i9991_2_lut_3_lut_4_lut_4_lut.init = 16'h8088;
    LUT4 i2_4_lut_adj_264 (.A(escape), .B(n31599), .C(n29647), .D(rx_data[6]), 
         .Z(n7_adj_186)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2_4_lut_adj_264.init = 16'h0004;
    LUT4 i22088_3_lut (.A(rx_data[5]), .B(rx_data[7]), .C(rx_data[3]), 
         .Z(n29647)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22088_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_265 (.A(n1473[4]), .B(\buffer[0] [0]), .C(n11_c), 
         .D(n14_c), .Z(n28592)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_265.init = 16'heca0;
    LUT4 reduce_or_462_i1_3_lut_4_lut (.A(n31522), .B(n13489), .C(\buffer[0] [7]), 
         .D(n1473[9]), .Z(n1578)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_462_i1_3_lut_4_lut.init = 16'hff80;
    PFUMX i38 (.BLUT(n25), .ALUT(n19), .C0(register_addr[0]), .Z(n28));
    LUT4 i1_4_lut_adj_266 (.A(n5833), .B(n13_adj_151), .C(n31500), .D(n1491), 
         .Z(n16767)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_266.init = 16'h8000;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_57)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 esc_data_2__bdd_4_lut (.A(esc_data[2]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[4]), .Z(n30733)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam esc_data_2__bdd_4_lut.init = 16'h4801;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_56)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_55)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_c)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_adj_267 (.A(\register[2] [3]), .B(n112), .C(n19331), 
         .D(n28899), .Z(n6002)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_267.init = 16'h333b;
    LUT4 i1_4_lut_adj_268 (.A(register_addr[1]), .B(n31505), .C(register_addr[0]), 
         .D(register_addr[2]), .Z(n112)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_268.init = 16'hfeff;
    LUT4 i2_3_lut_adj_269 (.A(register_addr[2]), .B(register_addr[3]), .C(n31523), 
         .Z(n28899)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_adj_269.init = 16'hfefe;
    LUT4 i22354_4_lut (.A(n31538), .B(n31589), .C(register_addr[2]), .D(n31590), 
         .Z(n27427)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i22354_4_lut.init = 16'h0111;
    LUT4 mux_1598_i24_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[23]), 
         .D(n224_adj_91[23]), .Z(n4094[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i25_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[24]), 
         .D(n224[24]), .Z(n3921[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i24_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[23]), 
         .D(n224[23]), .Z(n3921[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i23_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[22]), 
         .D(n224_adj_91[22]), .Z(n4094[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i22_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[21]), 
         .D(n224_adj_91[21]), .Z(n4094[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i20_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[19]), 
         .D(n224[19]), .Z(n3921[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i20_3_lut_4_lut.init = 16'hf780;
    PFUMX i21 (.BLUT(n12_adj_172), .ALUT(n6_adj_173), .C0(register_addr[0]), 
          .Z(n28826));
    LUT4 i1_2_lut_adj_270 (.A(register_addr[0]), .B(\control_reg[7]_adj_37 ), 
         .Z(n8653)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_270.init = 16'h4444;
    LUT4 mux_1598_i21_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[20]), 
         .D(n224_adj_91[20]), .Z(n4094[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i22322_4_lut (.A(n7_adj_125), .B(n29559), .C(n31551), .D(n1473[3]), 
         .Z(n13041)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i22322_4_lut.init = 16'h0544;
    LUT4 i22005_3_lut (.A(n1473[13]), .B(n1473[0]), .C(n1473[4]), .Z(n29559)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22005_3_lut.init = 16'hfefe;
    LUT4 mux_1598_i12_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[11]), 
         .D(n224_adj_91[11]), .Z(n4094[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i11_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[10]), 
         .D(n224_adj_91[10]), .Z(n4094[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i10_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[9]), 
         .D(n224_adj_91[9]), .Z(n4094[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1598_i9_3_lut_4_lut (.A(n31415), .B(n31422), .C(databus[8]), 
         .D(n224_adj_91[8]), .Z(n4094[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1598_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1553_i22_3_lut_4_lut (.A(n31414), .B(n31422), .C(databus[21]), 
         .D(n224[21]), .Z(n3921[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1553_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_271 (.A(n29423), .B(n31599), .C(escape), .D(n30735), 
         .Z(n29228)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_271.init = 16'hccc8;
    LUT4 reduce_or_468_i1_3_lut (.A(busy), .B(n1473[13]), .C(n1485), .Z(n1584)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_468_i1_3_lut.init = 16'hdcdc;
    LUT4 i470_2_lut (.A(n5833), .B(n1491), .Z(n1585)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i470_2_lut.init = 16'h4444;
    PFUMX i23003 (.BLUT(n31644), .ALUT(n31645), .C0(n1926), .Z(n31646));
    PFUMX i23001 (.BLUT(n31641), .ALUT(n31642), .C0(n1926), .Z(n31643));
    PFUMX i22999 (.BLUT(n31638), .ALUT(n31639), .C0(sendcount[0]), .Z(n31640));
    PFUMX i22997 (.BLUT(n31635), .ALUT(n31636), .C0(sendcount[0]), .Z(n31637));
    PFUMX i22995 (.BLUT(n31632), .ALUT(n31633), .C0(sendcount[0]), .Z(n31634));
    PFUMX i22993 (.BLUT(n31629), .ALUT(n31630), .C0(sendcount[0]), .Z(n31631));
    PFUMX i22991 (.BLUT(n31626), .ALUT(n31627), .C0(sendcount[0]), .Z(n31628));
    PFUMX i22989 (.BLUT(n31623), .ALUT(n31624), .C0(sendcount[0]), .Z(n31625));
    LUT4 i1_2_lut_adj_272 (.A(rx_data[5]), .B(rx_data[0]), .Z(n29423)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_272.init = 16'hbbbb;
    PFUMX i22987 (.BLUT(n31620), .ALUT(n31621), .C0(sendcount[0]), .Z(n31622));
    LUT4 i4451_3_lut (.A(n1473[16]), .B(n2746), .C(busy), .Z(n11216)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4451_3_lut.init = 16'hcece;
    PFUMX i22985 (.BLUT(n31617), .ALUT(n31618), .C0(sendcount[3]), .Z(n5833));
    LUT4 i5580_3_lut (.A(busy), .B(n1488), .C(n1473[16]), .Z(n12347)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5580_3_lut.init = 16'ha8a8;
    LUT4 i2_4_lut_adj_273 (.A(n38), .B(busy), .C(n30341), .D(n1488), 
         .Z(n28604)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_273.init = 16'hfbfa;
    PFUMX i22981 (.BLUT(n31611), .ALUT(n31612), .C0(sendcount[0]), .Z(n31613));
    PFUMX i22979 (.BLUT(n31608), .ALUT(n31609), .C0(n31450), .Z(n31610));
    \UARTTransmitter(baud_div=12)  uart_output (.n33389(n33389), .tx_data({tx_data}), 
            .send(send), .\state[3] (\state[3] ), .\state[1] (\state[1] ), 
            .\state[0] (\state[0] ), .n1155(n1155), .n73(n73), .n31500(n31500), 
            .busy(busy), .n31472(n31472), .\reset_count[7] (\reset_count[7] ), 
            .\reset_count[6] (\reset_count[6] ), .\reset_count[5] (\reset_count[5] ), 
            .n27249(n27249), .n11072(n11072), .debug_c_c(debug_c_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_c(debug_c_c), .n31500(n31500), 
            .rx_data({rx_data}), .n33389(n33389), .uart_rx_c(uart_rx_c), 
            .debug_c_7(debug_c_7), .n29423(n29423), .n29276(n29276), .n57(n57_adj_109), 
            .n31453(n31453), .n30735(n30735), .n31472(n31472), .n1501(n1473[4]), 
            .n1503(n1473[2]), .n13464(n13464), .n1505(n1473[0]), .escape(escape), 
            .n1502(n1473[3]), .n12481(n12481), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (n33389, tx_data, send, \state[3] , 
            \state[1] , \state[0] , n1155, n73, n31500, busy, n31472, 
            \reset_count[7] , \reset_count[6] , \reset_count[5] , n27249, 
            n11072, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    input n33389;
    input [7:0]tx_data;
    input send;
    input \state[3] ;
    input \state[1] ;
    input \state[0] ;
    input n1155;
    output n73;
    input n31500;
    output busy;
    input n31472;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n27249;
    output n11072;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n30445, n30317;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9450, n30769, n14986, n31187, n31597, n31186, n42, n29731, 
        n29732, n30316, n30315, n28968, n31314, n7, n10, n104, 
        n12, n28971, n40, n29733, n2;
    
    LUT4 state_1__bdd_4_lut_22673 (.A(state[1]), .B(state[0]), .C(state[3]), 
         .D(state[2]), .Z(n30445)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam state_1__bdd_4_lut_22673.init = 16'h0f7e;
    FD1S3IX state__i0 (.D(n30317), .CK(bclk), .CD(n33389), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9450), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(send), .Z(n30769)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h7ffe;
    LUT4 i71_4_lut_4_lut (.A(\state[3] ), .B(\state[1] ), .C(\state[0] ), 
         .D(n1155), .Z(n73)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i71_4_lut_4_lut.init = 16'h8001;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n30769), .B(state[2]), .C(n31500), .Z(n14986)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'hefef;
    FD1P3IX busy_34 (.D(n31597), .SP(n31187), .CD(n31472), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 n31186_bdd_2_lut (.A(n31186), .B(state[2]), .Z(n31187)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n31186_bdd_2_lut.init = 16'h2222;
    LUT4 send_bdd_4_lut (.A(send), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n31186)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)))) */ ;
    defparam send_bdd_4_lut.init = 16'hc002;
    LUT4 i1_2_lut (.A(state[1]), .B(state[0]), .Z(n42)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i22171_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n29731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22171_3_lut.init = 16'hcaca;
    LUT4 i22172_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n29732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22172_3_lut.init = 16'hcaca;
    LUT4 state_3__bdd_4_lut (.A(state[3]), .B(state[0]), .C(send), .D(state[1]), 
         .Z(n30316)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;
    defparam state_3__bdd_4_lut.init = 16'hb332;
    LUT4 state_3__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n30315)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_3__bdd_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[0]), .C(n31500), .Z(n28968)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 n2801_bdd_4_lut (.A(n31500), .B(state[3]), .C(n42), .D(state[2]), 
         .Z(n31314)) /* synthesis lut_function=(!((B (D)+!B !(C (D)))+!A)) */ ;
    defparam n2801_bdd_4_lut.init = 16'h2088;
    LUT4 i2_3_lut (.A(\reset_count[7] ), .B(\reset_count[6] ), .C(\reset_count[5] ), 
         .Z(n27249)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    FD1P3AX state__i3 (.D(n31314), .SP(n14986), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9450), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9450), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9450), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9450), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9450), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9450), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9450), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i13087_1_lut_rep_454 (.A(state[3]), .Z(n31597)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i13087_1_lut_rep_454.init = 16'h5555;
    LUT4 i1_4_lut (.A(n31500), .B(state[3]), .C(n12), .D(state[2]), 
         .Z(n28971)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam i1_4_lut.init = 16'h20a0;
    LUT4 i22_2_lut (.A(state[1]), .B(state[0]), .Z(n12)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i22_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_4_lut (.A(state[3]), .B(state[2]), .C(n42), .D(n31500), 
         .Z(n40)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut_4_lut.init = 16'h3400;
    PFUMX i22173 (.BLUT(n29731), .ALUT(n29732), .C0(state[1]), .Z(n29733));
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n29733), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15243_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15243_4_lut.init = 16'hfcee;
    FD1P3AX state__i2 (.D(n40), .SP(n14986), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n28971), .SP(n14986), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3JX tx_35 (.D(n104), .SP(n30445), .PD(n33389), .CK(bclk), .Q(n11072)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(send), .B(state[3]), .C(state[1]), .D(n28968), 
         .Z(n9450)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i3_4_lut.init = 16'h0200;
    PFUMX i22574 (.BLUT(n30316), .ALUT(n30315), .C0(state[2]), .Z(n30317));
    \ClockDividerP(factor=12)  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (bclk, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n8471, n27082, n27081;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27080, n27079, n27078, n27077, n27076, n27075, n27074, 
        n27073, n27072, n27071, n27070, n27069, n27068, n27067, 
        n55, n56, n4, n16803, n52, n44, n35, n54, n48, n36, 
        n46, n32;
    wire [31:0]n102;
    
    wire n50, n40, n27018, n27017, n27016, n27015, n27014, n27013, 
        n27012, n27011, n27010, n27009, n27008, n27007, n27006, 
        n27005, n27004, n27003;
    
    FD1S3AX clk_o_14 (.D(n8471), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D sub_2085_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27082), .S0(n8471));
    defparam sub_2085_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2085_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2085_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2085_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27081), .COUT(n27082));
    defparam sub_2085_add_2_32.INIT0 = 16'h5555;
    defparam sub_2085_add_2_32.INIT1 = 16'h5555;
    defparam sub_2085_add_2_32.INJECT1_0 = "NO";
    defparam sub_2085_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27080), .COUT(n27081));
    defparam sub_2085_add_2_30.INIT0 = 16'h5555;
    defparam sub_2085_add_2_30.INIT1 = 16'h5555;
    defparam sub_2085_add_2_30.INJECT1_0 = "NO";
    defparam sub_2085_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27079), .COUT(n27080));
    defparam sub_2085_add_2_28.INIT0 = 16'h5555;
    defparam sub_2085_add_2_28.INIT1 = 16'h5555;
    defparam sub_2085_add_2_28.INJECT1_0 = "NO";
    defparam sub_2085_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27078), .COUT(n27079));
    defparam sub_2085_add_2_26.INIT0 = 16'h5555;
    defparam sub_2085_add_2_26.INIT1 = 16'h5555;
    defparam sub_2085_add_2_26.INJECT1_0 = "NO";
    defparam sub_2085_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27077), .COUT(n27078));
    defparam sub_2085_add_2_24.INIT0 = 16'h5555;
    defparam sub_2085_add_2_24.INIT1 = 16'h5555;
    defparam sub_2085_add_2_24.INJECT1_0 = "NO";
    defparam sub_2085_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27076), .COUT(n27077));
    defparam sub_2085_add_2_22.INIT0 = 16'h5555;
    defparam sub_2085_add_2_22.INIT1 = 16'h5555;
    defparam sub_2085_add_2_22.INJECT1_0 = "NO";
    defparam sub_2085_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27075), .COUT(n27076));
    defparam sub_2085_add_2_20.INIT0 = 16'h5555;
    defparam sub_2085_add_2_20.INIT1 = 16'h5555;
    defparam sub_2085_add_2_20.INJECT1_0 = "NO";
    defparam sub_2085_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27074), .COUT(n27075));
    defparam sub_2085_add_2_18.INIT0 = 16'h5555;
    defparam sub_2085_add_2_18.INIT1 = 16'h5555;
    defparam sub_2085_add_2_18.INJECT1_0 = "NO";
    defparam sub_2085_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27073), .COUT(n27074));
    defparam sub_2085_add_2_16.INIT0 = 16'h5555;
    defparam sub_2085_add_2_16.INIT1 = 16'h5555;
    defparam sub_2085_add_2_16.INJECT1_0 = "NO";
    defparam sub_2085_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27072), .COUT(n27073));
    defparam sub_2085_add_2_14.INIT0 = 16'h5555;
    defparam sub_2085_add_2_14.INIT1 = 16'h5555;
    defparam sub_2085_add_2_14.INJECT1_0 = "NO";
    defparam sub_2085_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27071), .COUT(n27072));
    defparam sub_2085_add_2_12.INIT0 = 16'h5555;
    defparam sub_2085_add_2_12.INIT1 = 16'h5555;
    defparam sub_2085_add_2_12.INJECT1_0 = "NO";
    defparam sub_2085_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27070), .COUT(n27071));
    defparam sub_2085_add_2_10.INIT0 = 16'h5555;
    defparam sub_2085_add_2_10.INIT1 = 16'h5555;
    defparam sub_2085_add_2_10.INJECT1_0 = "NO";
    defparam sub_2085_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27069), .COUT(n27070));
    defparam sub_2085_add_2_8.INIT0 = 16'h5555;
    defparam sub_2085_add_2_8.INIT1 = 16'h5555;
    defparam sub_2085_add_2_8.INJECT1_0 = "NO";
    defparam sub_2085_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27068), .COUT(n27069));
    defparam sub_2085_add_2_6.INIT0 = 16'h5555;
    defparam sub_2085_add_2_6.INIT1 = 16'h5555;
    defparam sub_2085_add_2_6.INJECT1_0 = "NO";
    defparam sub_2085_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27067), .COUT(n27068));
    defparam sub_2085_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2085_add_2_4.INIT1 = 16'h5555;
    defparam sub_2085_add_2_4.INJECT1_0 = "NO";
    defparam sub_2085_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2085_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27067));
    defparam sub_2085_add_2_2.INIT0 = 16'h0000;
    defparam sub_2085_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2085_add_2_2.INJECT1_0 = "NO";
    defparam sub_2085_add_2_2.INJECT1_1 = "NO";
    LUT4 i22382_4_lut (.A(n55), .B(count[1]), .C(n56), .D(n4), .Z(n16803)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22382_4_lut.init = 16'h0400;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[3]), .B(count[0]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i6_2_lut.init = 16'heeee;
    FD1S3IX count_2678__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i0.GSR = "ENABLED";
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i11_2_lut.init = 16'heeee;
    FD1S3IX count_2678__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i1.GSR = "ENABLED";
    FD1S3IX count_2678__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i2.GSR = "ENABLED";
    FD1S3IX count_2678__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i3.GSR = "ENABLED";
    FD1S3IX count_2678__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i4.GSR = "ENABLED";
    FD1S3IX count_2678__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i5.GSR = "ENABLED";
    FD1S3IX count_2678__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i6.GSR = "ENABLED";
    FD1S3IX count_2678__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i7.GSR = "ENABLED";
    FD1S3IX count_2678__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i8.GSR = "ENABLED";
    FD1S3IX count_2678__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i9.GSR = "ENABLED";
    FD1S3IX count_2678__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i10.GSR = "ENABLED";
    FD1S3IX count_2678__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i11.GSR = "ENABLED";
    FD1S3IX count_2678__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i12.GSR = "ENABLED";
    FD1S3IX count_2678__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i13.GSR = "ENABLED";
    FD1S3IX count_2678__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i14.GSR = "ENABLED";
    FD1S3IX count_2678__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i15.GSR = "ENABLED";
    FD1S3IX count_2678__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i16.GSR = "ENABLED";
    FD1S3IX count_2678__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i17.GSR = "ENABLED";
    FD1S3IX count_2678__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i18.GSR = "ENABLED";
    FD1S3IX count_2678__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i19.GSR = "ENABLED";
    FD1S3IX count_2678__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i20.GSR = "ENABLED";
    FD1S3IX count_2678__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i21.GSR = "ENABLED";
    FD1S3IX count_2678__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i22.GSR = "ENABLED";
    FD1S3IX count_2678__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i23.GSR = "ENABLED";
    FD1S3IX count_2678__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i24.GSR = "ENABLED";
    FD1S3IX count_2678__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i25.GSR = "ENABLED";
    FD1S3IX count_2678__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i26.GSR = "ENABLED";
    FD1S3IX count_2678__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i27.GSR = "ENABLED";
    FD1S3IX count_2678__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i28.GSR = "ENABLED";
    FD1S3IX count_2678__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i29.GSR = "ENABLED";
    FD1S3IX count_2678__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i30.GSR = "ENABLED";
    FD1S3IX count_2678__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16803), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i31.GSR = "ENABLED";
    CCU2D count_2678_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27018), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_33.INIT1 = 16'h0000;
    defparam count_2678_add_4_33.INJECT1_0 = "NO";
    defparam count_2678_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27017), .COUT(n27018), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_31.INJECT1_0 = "NO";
    defparam count_2678_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27016), .COUT(n27017), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_29.INJECT1_0 = "NO";
    defparam count_2678_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27015), .COUT(n27016), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_27.INJECT1_0 = "NO";
    defparam count_2678_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27014), .COUT(n27015), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_25.INJECT1_0 = "NO";
    defparam count_2678_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27013), .COUT(n27014), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_23.INJECT1_0 = "NO";
    defparam count_2678_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27012), .COUT(n27013), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_21.INJECT1_0 = "NO";
    defparam count_2678_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27011), .COUT(n27012), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_19.INJECT1_0 = "NO";
    defparam count_2678_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27010), .COUT(n27011), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_17.INJECT1_0 = "NO";
    defparam count_2678_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27009), .COUT(n27010), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_15.INJECT1_0 = "NO";
    defparam count_2678_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27008), .COUT(n27009), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_13.INJECT1_0 = "NO";
    defparam count_2678_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27007), .COUT(n27008), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_11.INJECT1_0 = "NO";
    defparam count_2678_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27006), .COUT(n27007), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_9.INJECT1_0 = "NO";
    defparam count_2678_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27005), .COUT(n27006), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_7.INJECT1_0 = "NO";
    defparam count_2678_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27004), .COUT(n27005), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_5.INJECT1_0 = "NO";
    defparam count_2678_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27003), .COUT(n27004), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_3.INJECT1_0 = "NO";
    defparam count_2678_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27003), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_1.INIT0 = 16'hF000;
    defparam count_2678_add_4_1.INIT1 = 16'h0555;
    defparam count_2678_add_4_1.INJECT1_0 = "NO";
    defparam count_2678_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_c, n31500, rx_data, n33389, 
            uart_rx_c, debug_c_7, n29423, n29276, n57, n31453, n30735, 
            n31472, n1501, n1503, n13464, n1505, escape, n1502, 
            n12481, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31500;
    output [7:0]rx_data;
    input n33389;
    input uart_rx_c;
    output debug_c_7;
    input n29423;
    input n29276;
    output n57;
    output n31453;
    output n30735;
    input n31472;
    input n1501;
    input n1503;
    output n13464;
    input n1505;
    input escape;
    input n1502;
    output n12481;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n9398, n9400;
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n28512, baud_reset, n19, n31560, n31519, n31497, n31490, 
        n31568, n31562, n13568, n19_adj_32, n30709, n30708, n31403;
    wire [7:0]n78;
    
    wire n13559, n13, n9414, n31602, n9416, n31567, n29322, n9418, 
        n9420, n29383, n9422, n22200, n9424, n9426, n10238, bclk, 
        n29202, n16636, n30788, n9428, n9430, n9432, n9434, n9436, 
        n9438, n29371, n24508, n19_adj_33, n9440, n27, n28296, 
        n31513, n29392, n31518, n30734, n31566, n31498, n25, n27_adj_34, 
        n28398, n21, n23, n28050, n16637, n4, n4_adj_35, n51, 
        n47;
    
    FD1P3AX rdata_i0_i0 (.D(n9398), .SP(n31500), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n9400), .SP(n31500), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n28512), .CK(debug_c_c), .CD(n33389), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n19), .CK(debug_c_c), .PD(n33389), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_354_4_lut (.A(state[4]), .B(state[3]), .C(n31560), 
         .D(n31519), .Z(n31497)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_354_4_lut.init = 16'heaff;
    LUT4 i1_2_lut_rep_347_4_lut (.A(state[4]), .B(state[3]), .C(n31560), 
         .D(state[5]), .Z(n31490)) /* synthesis lut_function=(!(A (D)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_347_4_lut.init = 16'h00ea;
    LUT4 i2_3_lut_4_lut (.A(n31568), .B(n31562), .C(state[0]), .D(state[5]), 
         .Z(n13568)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_4_lut_adj_57 (.A(state[0]), .B(n31562), .C(state[5]), 
         .D(n31568), .Z(n19_adj_32)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_4_lut_adj_57.init = 16'hffef;
    LUT4 n30709_bdd_4_lut (.A(n30709), .B(state[5]), .C(n30708), .D(state[0]), 
         .Z(n31403)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam n30709_bdd_4_lut.init = 16'hf022;
    LUT4 i1_4_lut (.A(n78[1]), .B(rdata[1]), .C(n13559), .D(n13), .Z(n9414)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i4410_4_lut (.A(uart_rx_c), .B(rdata[1]), .C(n31568), .D(n31602), 
         .Z(n78[1])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4410_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_58 (.A(n78[2]), .B(rdata[2]), .C(n13559), .D(n13), 
         .Z(n9416)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_58.init = 16'heca0;
    LUT4 i4408_4_lut (.A(uart_rx_c), .B(rdata[2]), .C(n31567), .D(n29322), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4408_4_lut.init = 16'hccca;
    LUT4 i1_2_lut (.A(state[3]), .B(state[2]), .Z(n29322)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_59 (.A(n78[3]), .B(rdata[3]), .C(n13559), .D(n13), 
         .Z(n9418)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_59.init = 16'heca0;
    LUT4 i4406_4_lut (.A(uart_rx_c), .B(rdata[3]), .C(n31602), .D(n29322), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4406_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_60 (.A(n78[4]), .B(rdata[4]), .C(n13559), .D(n13), 
         .Z(n9420)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_60.init = 16'heca0;
    LUT4 i4404_4_lut (.A(uart_rx_c), .B(rdata[4]), .C(state[2]), .D(n29383), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4404_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_61 (.A(n78[5]), .B(rdata[5]), .C(n13559), .D(n13), 
         .Z(n9422)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_61.init = 16'heca0;
    LUT4 i4402_4_lut (.A(uart_rx_c), .B(rdata[5]), .C(state[2]), .D(n22200), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4402_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_62 (.A(n78[6]), .B(rdata[6]), .C(n13559), .D(n13), 
         .Z(n9424)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_62.init = 16'heca0;
    LUT4 i4400_4_lut (.A(uart_rx_c), .B(rdata[6]), .C(state[2]), .D(n29383), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4400_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_63 (.A(n78[7]), .B(rdata[7]), .C(n13559), .D(n13), 
         .Z(n9426)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_63.init = 16'heca0;
    LUT4 i1_4_lut_4_lut (.A(state[4]), .B(n10238), .C(bclk), .D(n31490), 
         .Z(n29202)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h6a00;
    LUT4 i9864_3_lut_3_lut (.A(state[4]), .B(n10238), .C(bclk), .Z(n16636)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i9864_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i4398_4_lut (.A(rdata[7]), .B(uart_rx_c), .C(state[2]), .D(n22200), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4398_4_lut.init = 16'hcaaa;
    LUT4 state_3__bdd_4_lut (.A(state[3]), .B(bclk), .C(state[2]), .D(state[1]), 
         .Z(n30788)) /* synthesis lut_function=(A (B+!(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam state_3__bdd_4_lut.init = 16'h9aaa;
    LUT4 i1_4_lut_adj_64 (.A(rdata[1]), .B(rx_data[1]), .C(n13568), .D(n19_adj_32), 
         .Z(n9428)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_64.init = 16'heca0;
    LUT4 i1_4_lut_adj_65 (.A(rdata[2]), .B(rx_data[2]), .C(n13568), .D(n19_adj_32), 
         .Z(n9430)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_65.init = 16'heca0;
    LUT4 i1_4_lut_adj_66 (.A(rdata[3]), .B(rx_data[3]), .C(n13568), .D(n19_adj_32), 
         .Z(n9432)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_66.init = 16'heca0;
    LUT4 i1_4_lut_adj_67 (.A(rdata[4]), .B(rx_data[4]), .C(n13568), .D(n19_adj_32), 
         .Z(n9434)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_67.init = 16'heca0;
    LUT4 i1_4_lut_adj_68 (.A(rdata[5]), .B(rx_data[5]), .C(n13568), .D(n19_adj_32), 
         .Z(n9436)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_68.init = 16'heca0;
    LUT4 i1_4_lut_adj_69 (.A(rdata[6]), .B(rx_data[6]), .C(n13568), .D(n19_adj_32), 
         .Z(n9438)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_69.init = 16'heca0;
    LUT4 i22422_4_lut (.A(debug_c_7), .B(n29371), .C(uart_rx_c), .D(n24508), 
         .Z(n19_adj_33)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i22422_4_lut.init = 16'ha8ec;
    LUT4 i1_4_lut_adj_70 (.A(rdata[7]), .B(rx_data[7]), .C(n13568), .D(n19_adj_32), 
         .Z(n9440)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_70.init = 16'heca0;
    LUT4 i43_4_lut (.A(state[5]), .B(n30788), .C(state[0]), .D(n27), 
         .Z(n28296)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i43_4_lut.init = 16'hc5c0;
    LUT4 i2_3_lut_4_lut_adj_71 (.A(n31513), .B(n29423), .C(rx_data[3]), 
         .D(n29276), .Z(n57)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut_adj_71.init = 16'h1000;
    LUT4 i2_3_lut_rep_310_4_lut (.A(n31513), .B(n29423), .C(rx_data[1]), 
         .D(n29392), .Z(n31453)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_310_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut (.A(state[5]), .B(n31518), .C(state[0]), .D(bclk), 
         .Z(n28512)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut.init = 16'hf400;
    LUT4 n30734_bdd_2_lut_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(n30734), 
         .Z(n30735)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam n30734_bdd_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_370_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(rx_data[2]), 
         .Z(n31513)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_370_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_4_lut (.A(uart_rx_c), .B(n31519), .C(state[3]), 
         .D(n31518), .Z(n27)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A ((C (D))+!B)) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hf131;
    FD1S3IX drdy_51 (.D(n19_adj_33), .CK(debug_c_c), .CD(n31472), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_417 (.A(state[1]), .B(state[2]), .Z(n31560)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_417.init = 16'h8888;
    LUT4 i1_3_lut_rep_375_4_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .D(state[4]), .Z(n31518)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut_rep_375_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_419 (.A(state[1]), .B(state[4]), .Z(n31562)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_419.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(n31566), 
         .D(n31568), .Z(n29371)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21903_2_lut_rep_355_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(uart_rx_c), 
         .D(n31568), .Z(n31498)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21903_2_lut_rep_355_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_72 (.A(state[1]), .B(state[4]), .C(n31568), 
         .D(state[0]), .Z(n24508)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut_adj_72.init = 16'hfffe;
    PFUMX i40 (.BLUT(n25), .ALUT(n27_adj_34), .C0(state[0]), .Z(n28398));
    LUT4 i14720_2_lut_rep_423 (.A(state[0]), .B(state[5]), .Z(n31566)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14720_2_lut_rep_423.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13559)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_424 (.A(state[1]), .B(bclk), .Z(n31567)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_rep_424.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_73 (.A(state[1]), .B(bclk), .C(state[3]), 
         .Z(n29383)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_3_lut_adj_73.init = 16'hbfbf;
    LUT4 i2_2_lut_rep_425 (.A(state[3]), .B(state[2]), .Z(n31568)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_2_lut_rep_425.init = 16'heeee;
    LUT4 i1_2_lut_rep_376_3_lut_4_lut (.A(state[3]), .B(state[2]), .C(state[4]), 
         .D(state[1]), .Z(n31519)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_376_3_lut_4_lut.init = 16'hfffe;
    LUT4 state_1__bdd_2_lut (.A(state[1]), .B(bclk), .Z(n30708)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam state_1__bdd_2_lut.init = 16'h9999;
    PFUMX i36 (.BLUT(n21), .ALUT(n23), .C0(state[5]), .Z(n28050));
    PFUMX i9865 (.BLUT(n29202), .ALUT(n16636), .C0(state[0]), .Z(n16637));
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(n31518), .C(n31519), .D(uart_rx_c), 
         .Z(n30709)) /* synthesis lut_function=(A (B+!(C))+!A !(C+(D))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8a8f;
    LUT4 i41_4_lut_3_lut (.A(bclk), .B(state[1]), .C(state[2]), .Z(n27_adj_34)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i41_4_lut_3_lut.init = 16'hb4b4;
    LUT4 i1_4_lut_adj_74 (.A(rdata[0]), .B(rx_data[0]), .C(n13568), .D(n19_adj_32), 
         .Z(n9400)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_74.init = 16'heca0;
    FD1P3AX rdata_i0_i1 (.D(n9414), .SP(n31500), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n9416), .SP(n31500), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n9418), .SP(n31500), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n9420), .SP(n31500), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n9422), .SP(n31500), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n9424), .SP(n31500), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n9426), .SP(n31500), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n9428), .SP(n31500), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n9430), .SP(n31500), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n9432), .SP(n31500), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n9434), .SP(n31500), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n9436), .SP(n31500), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n9438), .SP(n31500), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n9440), .SP(n31500), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n31403), .CK(debug_c_c), .CD(n31472), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n28398), .CK(debug_c_c), .CD(n31472), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n28296), .CK(debug_c_c), .CD(n31472), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n16637), .CK(debug_c_c), .CD(n31472), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n28050), .CK(debug_c_c), .CD(n31472), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_75 (.A(state[5]), .B(n31498), .C(state[2]), .D(n31497), 
         .Z(n25)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_75.init = 16'h5111;
    LUT4 i15064_2_lut_rep_459 (.A(bclk), .B(state[1]), .Z(n31602)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15064_2_lut_rep_459.init = 16'h8888;
    LUT4 i15468_2_lut_3_lut (.A(bclk), .B(state[1]), .C(state[3]), .Z(n22200)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15468_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_4_lut (.A(bclk), .B(n4), .C(state[0]), .D(n31518), .Z(n21)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'h4840;
    LUT4 i1_2_lut_adj_76 (.A(state[4]), .B(n10238), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_76.init = 16'h8888;
    LUT4 i38_4_lut (.A(n31498), .B(n10238), .C(state[0]), .D(n4_adj_35), 
         .Z(n23)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i38_4_lut.init = 16'hf535;
    LUT4 i1_2_lut_adj_77 (.A(state[4]), .B(bclk), .Z(n4_adj_35)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_77.init = 16'hdddd;
    LUT4 i22426_4_lut (.A(baud_reset), .B(n29371), .C(uart_rx_c), .D(n24508), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i22426_4_lut.init = 16'ha8ec;
    LUT4 i3447_4_lut (.A(state[3]), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(n10238)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3447_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_78 (.A(n78[0]), .B(rdata[0]), .C(n13559), .D(n13), 
         .Z(n9398)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_78.init = 16'heca0;
    LUT4 i4453_4_lut (.A(uart_rx_c), .B(rdata[0]), .C(n31568), .D(n31567), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4453_4_lut.init = 16'hccca;
    LUT4 i2_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut.init = 16'hefef;
    LUT4 rx_data_1__bdd_4_lut (.A(rx_data[1]), .B(rx_data[3]), .C(rx_data[4]), 
         .D(rx_data[2]), .Z(n30734)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C (D)))+!A (B+(C+(D)))) */ ;
    defparam rx_data_1__bdd_4_lut.init = 16'hdf7e;
    LUT4 i1_4_lut_adj_79 (.A(n1501), .B(debug_c_7), .C(n1503), .D(n51), 
         .Z(n13464)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_79.init = 16'heeea;
    LUT4 i47_4_lut (.A(n31453), .B(n1505), .C(n47), .D(n57), .Z(n51)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i47_4_lut.init = 16'h4f45;
    LUT4 i1_2_lut_adj_80 (.A(escape), .B(n1502), .Z(n47)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_80.init = 16'hbbbb;
    LUT4 i1_3_lut (.A(debug_c_7), .B(n1503), .C(n1502), .Z(n12481)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i1_3_lut.init = 16'h5454;
    LUT4 i1_2_lut_adj_81 (.A(rx_data[4]), .B(rx_data[3]), .Z(n29392)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_81.init = 16'heeee;
    \ClockDividerP(factor=12)_U0  baud_gen (.GND_net(GND_net), .baud_reset(baud_reset), 
            .bclk(bclk), .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (GND_net, baud_reset, bclk, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input baud_reset;
    output bclk;
    input debug_c_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26986;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n26985, n26984, n26983, n26982, n26981, n26980, n26979, 
        n26978, n26977, n26976, n26975, n26974, n26973, n26972, 
        n26971, n57, n55, n56, n2962, n54, n46, n29623, n50, 
        n38, n52, n42, n48, n34, n8436, n27098, n27097, n27096, 
        n27095, n27094, n27093, n27092, n27091, n27090, n27089, 
        n27088, n27087, n27086, n27085, n27084, n27083;
    
    CCU2D count_2677_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26986), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_33.INIT1 = 16'h0000;
    defparam count_2677_add_4_33.INJECT1_0 = "NO";
    defparam count_2677_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26985), .COUT(n26986), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_31.INJECT1_0 = "NO";
    defparam count_2677_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26984), .COUT(n26985), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_29.INJECT1_0 = "NO";
    defparam count_2677_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26983), .COUT(n26984), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_27.INJECT1_0 = "NO";
    defparam count_2677_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26982), .COUT(n26983), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_25.INJECT1_0 = "NO";
    defparam count_2677_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26981), .COUT(n26982), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_23.INJECT1_0 = "NO";
    defparam count_2677_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26980), .COUT(n26981), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_21.INJECT1_0 = "NO";
    defparam count_2677_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26979), .COUT(n26980), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_19.INJECT1_0 = "NO";
    defparam count_2677_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26978), .COUT(n26979), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_17.INJECT1_0 = "NO";
    defparam count_2677_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26977), .COUT(n26978), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_15.INJECT1_0 = "NO";
    defparam count_2677_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26976), .COUT(n26977), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_13.INJECT1_0 = "NO";
    defparam count_2677_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26975), .COUT(n26976), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_11.INJECT1_0 = "NO";
    defparam count_2677_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26974), .COUT(n26975), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_9.INJECT1_0 = "NO";
    defparam count_2677_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26973), .COUT(n26974), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_7.INJECT1_0 = "NO";
    defparam count_2677_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26972), .COUT(n26973), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_5.INJECT1_0 = "NO";
    defparam count_2677_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26971), .COUT(n26972), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_3.INJECT1_0 = "NO";
    defparam count_2677_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26971), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677_add_4_1.INIT0 = 16'hF000;
    defparam count_2677_add_4_1.INIT1 = 16'h0555;
    defparam count_2677_add_4_1.INJECT1_0 = "NO";
    defparam count_2677_add_4_1.INJECT1_1 = "NO";
    LUT4 i1112_4_lut (.A(n57), .B(baud_reset), .C(n55), .D(n56), .Z(n2962)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i1112_4_lut.init = 16'hcccd;
    LUT4 i27_4_lut (.A(count[31]), .B(n54), .C(n46), .D(n29623), .Z(n57)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i27_4_lut.init = 16'hfeff;
    LUT4 i25_4_lut (.A(count[24]), .B(n50), .C(n38), .D(count[4]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(count[5]), .B(n52), .C(n42), .D(count[6]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(count[16]), .B(n48), .C(n34), .D(count[11]), 
         .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(count[28]), .B(count[2]), .C(count[18]), .D(count[8]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i22064_3_lut (.A(count[3]), .B(count[0]), .C(count[1]), .Z(n29623)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22064_3_lut.init = 16'h8080;
    LUT4 i18_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[21]), .B(count[25]), .Z(n34)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i4_2_lut.init = 16'heeee;
    FD1S3IX clk_o_14 (.D(n8436), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    LUT4 i20_4_lut (.A(count[7]), .B(count[19]), .C(count[14]), .D(count[22]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(count[27]), .B(count[30]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(count[15]), .B(count[29]), .C(count[23]), .D(count[13]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i12_2_lut (.A(count[10]), .B(count[20]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_2_lut.init = 16'heeee;
    FD1S3IX count_2677__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2962), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i0.GSR = "ENABLED";
    CCU2D sub_2083_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27098), .S0(n8436));
    defparam sub_2083_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2083_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2083_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2083_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27097), .COUT(n27098));
    defparam sub_2083_add_2_32.INIT0 = 16'h5555;
    defparam sub_2083_add_2_32.INIT1 = 16'h5555;
    defparam sub_2083_add_2_32.INJECT1_0 = "NO";
    defparam sub_2083_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27096), .COUT(n27097));
    defparam sub_2083_add_2_30.INIT0 = 16'h5555;
    defparam sub_2083_add_2_30.INIT1 = 16'h5555;
    defparam sub_2083_add_2_30.INJECT1_0 = "NO";
    defparam sub_2083_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27095), .COUT(n27096));
    defparam sub_2083_add_2_28.INIT0 = 16'h5555;
    defparam sub_2083_add_2_28.INIT1 = 16'h5555;
    defparam sub_2083_add_2_28.INJECT1_0 = "NO";
    defparam sub_2083_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27094), .COUT(n27095));
    defparam sub_2083_add_2_26.INIT0 = 16'h5555;
    defparam sub_2083_add_2_26.INIT1 = 16'h5555;
    defparam sub_2083_add_2_26.INJECT1_0 = "NO";
    defparam sub_2083_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27093), .COUT(n27094));
    defparam sub_2083_add_2_24.INIT0 = 16'h5555;
    defparam sub_2083_add_2_24.INIT1 = 16'h5555;
    defparam sub_2083_add_2_24.INJECT1_0 = "NO";
    defparam sub_2083_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27092), .COUT(n27093));
    defparam sub_2083_add_2_22.INIT0 = 16'h5555;
    defparam sub_2083_add_2_22.INIT1 = 16'h5555;
    defparam sub_2083_add_2_22.INJECT1_0 = "NO";
    defparam sub_2083_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27091), .COUT(n27092));
    defparam sub_2083_add_2_20.INIT0 = 16'h5555;
    defparam sub_2083_add_2_20.INIT1 = 16'h5555;
    defparam sub_2083_add_2_20.INJECT1_0 = "NO";
    defparam sub_2083_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27090), .COUT(n27091));
    defparam sub_2083_add_2_18.INIT0 = 16'h5555;
    defparam sub_2083_add_2_18.INIT1 = 16'h5555;
    defparam sub_2083_add_2_18.INJECT1_0 = "NO";
    defparam sub_2083_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27089), .COUT(n27090));
    defparam sub_2083_add_2_16.INIT0 = 16'h5555;
    defparam sub_2083_add_2_16.INIT1 = 16'h5555;
    defparam sub_2083_add_2_16.INJECT1_0 = "NO";
    defparam sub_2083_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27088), .COUT(n27089));
    defparam sub_2083_add_2_14.INIT0 = 16'h5555;
    defparam sub_2083_add_2_14.INIT1 = 16'h5555;
    defparam sub_2083_add_2_14.INJECT1_0 = "NO";
    defparam sub_2083_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27087), .COUT(n27088));
    defparam sub_2083_add_2_12.INIT0 = 16'h5555;
    defparam sub_2083_add_2_12.INIT1 = 16'h5555;
    defparam sub_2083_add_2_12.INJECT1_0 = "NO";
    defparam sub_2083_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27086), .COUT(n27087));
    defparam sub_2083_add_2_10.INIT0 = 16'h5555;
    defparam sub_2083_add_2_10.INIT1 = 16'h5555;
    defparam sub_2083_add_2_10.INJECT1_0 = "NO";
    defparam sub_2083_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27085), .COUT(n27086));
    defparam sub_2083_add_2_8.INIT0 = 16'h5555;
    defparam sub_2083_add_2_8.INIT1 = 16'h5555;
    defparam sub_2083_add_2_8.INJECT1_0 = "NO";
    defparam sub_2083_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27084), .COUT(n27085));
    defparam sub_2083_add_2_6.INIT0 = 16'h5555;
    defparam sub_2083_add_2_6.INIT1 = 16'h5555;
    defparam sub_2083_add_2_6.INJECT1_0 = "NO";
    defparam sub_2083_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27083), .COUT(n27084));
    defparam sub_2083_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2083_add_2_4.INIT1 = 16'h5555;
    defparam sub_2083_add_2_4.INJECT1_0 = "NO";
    defparam sub_2083_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2083_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27083));
    defparam sub_2083_add_2_2.INIT0 = 16'h0000;
    defparam sub_2083_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2083_add_2_2.INJECT1_0 = "NO";
    defparam sub_2083_add_2_2.INJECT1_1 = "NO";
    FD1S3IX count_2677__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2962), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i1.GSR = "ENABLED";
    FD1S3IX count_2677__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2962), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i2.GSR = "ENABLED";
    FD1S3IX count_2677__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2962), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i3.GSR = "ENABLED";
    FD1S3IX count_2677__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2962), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i4.GSR = "ENABLED";
    FD1S3IX count_2677__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2962), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i5.GSR = "ENABLED";
    FD1S3IX count_2677__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2962), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i6.GSR = "ENABLED";
    FD1S3IX count_2677__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2962), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i7.GSR = "ENABLED";
    FD1S3IX count_2677__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2962), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i8.GSR = "ENABLED";
    FD1S3IX count_2677__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2962), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i9.GSR = "ENABLED";
    FD1S3IX count_2677__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i10.GSR = "ENABLED";
    FD1S3IX count_2677__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i11.GSR = "ENABLED";
    FD1S3IX count_2677__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i12.GSR = "ENABLED";
    FD1S3IX count_2677__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i13.GSR = "ENABLED";
    FD1S3IX count_2677__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i14.GSR = "ENABLED";
    FD1S3IX count_2677__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i15.GSR = "ENABLED";
    FD1S3IX count_2677__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i16.GSR = "ENABLED";
    FD1S3IX count_2677__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i17.GSR = "ENABLED";
    FD1S3IX count_2677__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i18.GSR = "ENABLED";
    FD1S3IX count_2677__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i19.GSR = "ENABLED";
    FD1S3IX count_2677__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i20.GSR = "ENABLED";
    FD1S3IX count_2677__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i21.GSR = "ENABLED";
    FD1S3IX count_2677__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i22.GSR = "ENABLED";
    FD1S3IX count_2677__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i23.GSR = "ENABLED";
    FD1S3IX count_2677__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i24.GSR = "ENABLED";
    FD1S3IX count_2677__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i25.GSR = "ENABLED";
    FD1S3IX count_2677__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i26.GSR = "ENABLED";
    FD1S3IX count_2677__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i27.GSR = "ENABLED";
    FD1S3IX count_2677__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i28.GSR = "ENABLED";
    FD1S3IX count_2677__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i29.GSR = "ENABLED";
    FD1S3IX count_2677__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i30.GSR = "ENABLED";
    FD1S3IX count_2677__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2962), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2677__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (\register[2] , GND_net, force_pause, debug_c_c, 
            n31511, \databus[1] , n9483, read_size, n14453, n31449, 
            prev_clk_1Hz, clk_1Hz, \register[0][2] , \select[1] , read_value, 
            n29068, rw, n46, n29292, n31477, n29293, n29294, n30305, 
            n30303, \reset_count[14] , n22483, xbee_pause_c, \register_addr[1] , 
            \register_addr[0] , n29169, n9537, n6002, n29065, n29055, 
            n29052, n16764, n27427, n29064, n16763, n29062, n29049, 
            n29051, n29053, n29066, n29056, n29067, n29070, n29071, 
            n29069, n6005, n29057, n29058, n29063, n29059, n29061, 
            n29054, n29050, n29048, n29060, n29047, n29788, n2875) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[2] ;
    input GND_net;
    output force_pause;
    input debug_c_c;
    input n31511;
    input \databus[1] ;
    input n9483;
    output [2:0]read_size;
    output n14453;
    input n31449;
    output prev_clk_1Hz;
    output clk_1Hz;
    output \register[0][2] ;
    input \select[1] ;
    output [31:0]read_value;
    input n29068;
    input rw;
    output n46;
    input n29292;
    input n31477;
    input n29293;
    input n29294;
    input n30305;
    input n30303;
    input \reset_count[14] ;
    input n22483;
    input xbee_pause_c;
    input \register_addr[1] ;
    input \register_addr[0] ;
    output n29169;
    input n9537;
    input n6002;
    input n29065;
    input n29055;
    input n29052;
    input n16764;
    input n27427;
    input n29064;
    input n16763;
    input n29062;
    input n29049;
    input n29051;
    input n29053;
    input n29066;
    input n29056;
    input n29067;
    input n29070;
    input n29071;
    input n29069;
    input n6005;
    input n29057;
    input n29058;
    input n29063;
    input n29059;
    input n29061;
    input n29054;
    input n29050;
    input n29048;
    input n29060;
    input n29047;
    output n29788;
    input n2875;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26724;
    wire [31:0]n100;
    
    wire n26725, n26723, n26722, n26721, n27236, n26720, n179, 
        prev_select, n26719, n26718, n26717, n26716, n26715, n31591, 
        n26730, n26729, n26728, n26727, n26726;
    
    CCU2D add_135_21 (.A0(\register[2] [19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26724), .COUT(n26725), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_21.INIT0 = 16'h5aaa;
    defparam add_135_21.INIT1 = 16'h5aaa;
    defparam add_135_21.INJECT1_0 = "NO";
    defparam add_135_21.INJECT1_1 = "NO";
    CCU2D add_135_19 (.A0(\register[2] [17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26723), .COUT(n26724), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_19.INIT0 = 16'h5aaa;
    defparam add_135_19.INIT1 = 16'h5aaa;
    defparam add_135_19.INJECT1_0 = "NO";
    defparam add_135_19.INJECT1_1 = "NO";
    CCU2D add_135_17 (.A0(\register[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26722), .COUT(n26723), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_17.INIT0 = 16'h5aaa;
    defparam add_135_17.INIT1 = 16'h5aaa;
    defparam add_135_17.INJECT1_0 = "NO";
    defparam add_135_17.INJECT1_1 = "NO";
    CCU2D add_135_15 (.A0(\register[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26721), .COUT(n26722), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_15.INIT0 = 16'h5aaa;
    defparam add_135_15.INIT1 = 16'h5aaa;
    defparam add_135_15.INJECT1_0 = "NO";
    defparam add_135_15.INJECT1_1 = "NO";
    FD1P3IX force_pause_152 (.D(\databus[1] ), .SP(n27236), .CD(n31511), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam force_pause_152.GSR = "ENABLED";
    CCU2D add_135_13 (.A0(\register[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26720), .COUT(n26721), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_13.INIT0 = 16'h5aaa;
    defparam add_135_13.INIT1 = 16'h5aaa;
    defparam add_135_13.INJECT1_0 = "NO";
    defparam add_135_13.INJECT1_1 = "NO";
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n9483), .CD(n31511), 
            .CK(debug_c_c), .Q(\register[2] [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n9483), .CD(n31511), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n31449), .SP(n14453), .CK(debug_c_c), 
            .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_150 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam prev_clk_1Hz_150.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_151 (.D(n179), .CK(debug_c_c), .Q(\register[0][2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam xbee_pause_latched_151.GSR = "ENABLED";
    FD1S3AX prev_select_149 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam prev_select_149.GSR = "ENABLED";
    CCU2D add_135_11 (.A0(\register[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26719), .COUT(n26720), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_11.INIT0 = 16'h5aaa;
    defparam add_135_11.INIT1 = 16'h5aaa;
    defparam add_135_11.INJECT1_0 = "NO";
    defparam add_135_11.INJECT1_1 = "NO";
    CCU2D add_135_9 (.A0(\register[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26718), .COUT(n26719), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_9.INIT0 = 16'h5aaa;
    defparam add_135_9.INIT1 = 16'h5aaa;
    defparam add_135_9.INJECT1_0 = "NO";
    defparam add_135_9.INJECT1_1 = "NO";
    CCU2D add_135_7 (.A0(\register[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26717), .COUT(n26718), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_7.INIT0 = 16'h5aaa;
    defparam add_135_7.INIT1 = 16'h5aaa;
    defparam add_135_7.INJECT1_0 = "NO";
    defparam add_135_7.INJECT1_1 = "NO";
    CCU2D add_135_5 (.A0(\register[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26716), .COUT(n26717), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_5.INIT0 = 16'h5aaa;
    defparam add_135_5.INIT1 = 16'h5aaa;
    defparam add_135_5.INJECT1_0 = "NO";
    defparam add_135_5.INJECT1_1 = "NO";
    CCU2D add_135_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26715), .COUT(n26716), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_3.INIT0 = 16'h5aaa;
    defparam add_135_3.INIT1 = 16'h5aaa;
    defparam add_135_3.INJECT1_0 = "NO";
    defparam add_135_3.INJECT1_1 = "NO";
    CCU2D add_135_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26715), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_1.INIT0 = 16'hF000;
    defparam add_135_1.INIT1 = 16'h5555;
    defparam add_135_1.INJECT1_0 = "NO";
    defparam add_135_1.INJECT1_1 = "NO";
    FD1P3AX read_value__i28 (.D(n29068), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i28.GSR = "ENABLED";
    LUT4 i14_2_lut (.A(\select[1] ), .B(rw), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(36[19:32])
    defparam i14_2_lut.init = 16'h8888;
    FD1P3AX read_value__i29 (.D(n29292), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i29.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n31511), .B(rw), .C(n31591), .D(n31477), .Z(n27236)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam i2_4_lut.init = 16'h0032;
    FD1P3AX read_value__i30 (.D(n29293), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n29294), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i2 (.D(n30305), .SP(n14453), .CK(debug_c_c), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3AX read_value__i1 (.D(n30303), .SP(n14453), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i118_2_lut_rep_448 (.A(prev_select), .B(\select[1] ), .Z(n31591)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(60[9:30])
    defparam i118_2_lut_rep_448.init = 16'h4444;
    LUT4 i964_2_lut_2_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(\reset_count[14] ), .D(n22483), .Z(n14453)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(60[9:30])
    defparam i964_2_lut_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i115_1_lut (.A(xbee_pause_c), .Z(n179)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(52[26:39])
    defparam i115_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n29169)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    FD1P3IX read_value__i3 (.D(n6002), .SP(n14453), .CD(n9537), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29065), .SP(n14453), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29055), .SP(n14453), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29052), .SP(n14453), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_size_i0_i1 (.D(n27427), .SP(n14453), .CD(n16764), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29064), .SP(n14453), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n31477), .SP(n14453), .CD(n16763), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29062), .SP(n14453), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29049), .SP(n14453), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29051), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29053), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29066), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29056), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29067), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29070), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29071), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29069), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n6005), .SP(n14453), .CD(n9537), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29057), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29058), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29063), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29059), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29061), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29054), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29050), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i24.GSR = "ENABLED";
    CCU2D add_135_33 (.A0(\register[2] [31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26730), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_33.INIT0 = 16'h5aaa;
    defparam add_135_33.INIT1 = 16'h0000;
    defparam add_135_33.INJECT1_0 = "NO";
    defparam add_135_33.INJECT1_1 = "NO";
    CCU2D add_135_31 (.A0(\register[2] [29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26729), .COUT(n26730), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_31.INIT0 = 16'h5aaa;
    defparam add_135_31.INIT1 = 16'h5aaa;
    defparam add_135_31.INJECT1_0 = "NO";
    defparam add_135_31.INJECT1_1 = "NO";
    FD1P3AX read_value__i25 (.D(n29048), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i25.GSR = "ENABLED";
    CCU2D add_135_29 (.A0(\register[2] [27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26728), .COUT(n26729), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_29.INIT0 = 16'h5aaa;
    defparam add_135_29.INIT1 = 16'h5aaa;
    defparam add_135_29.INJECT1_0 = "NO";
    defparam add_135_29.INJECT1_1 = "NO";
    CCU2D add_135_27 (.A0(\register[2] [25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26727), .COUT(n26728), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_27.INIT0 = 16'h5aaa;
    defparam add_135_27.INIT1 = 16'h5aaa;
    defparam add_135_27.INJECT1_0 = "NO";
    defparam add_135_27.INJECT1_1 = "NO";
    CCU2D add_135_25 (.A0(\register[2] [23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26726), .COUT(n26727), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_25.INIT0 = 16'h5aaa;
    defparam add_135_25.INIT1 = 16'h5aaa;
    defparam add_135_25.INJECT1_0 = "NO";
    defparam add_135_25.INJECT1_1 = "NO";
    FD1P3AX read_value__i26 (.D(n29060), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i26.GSR = "ENABLED";
    CCU2D add_135_23 (.A0(\register[2] [21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26725), .COUT(n26726), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_23.INIT0 = 16'h5aaa;
    defparam add_135_23.INIT1 = 16'h5aaa;
    defparam add_135_23.INJECT1_0 = "NO";
    defparam add_135_23.INJECT1_1 = "NO";
    FD1P3AX read_value__i27 (.D(n29047), .SP(n14453), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i27.GSR = "ENABLED";
    \ClockDividerP(factor=12000000)  uptime_div (.GND_net(GND_net), .clk_1Hz(clk_1Hz), 
            .debug_c_c(debug_c_c), .n31511(n31511), .n29788(n29788), .n2875(n2875)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(105[28] 107[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (GND_net, clk_1Hz, debug_c_c, 
            n31511, n29788, n2875) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output clk_1Hz;
    input debug_c_c;
    input n31511;
    output n29788;
    input n2875;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27180, n7985, n27179;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27178, n27177, n27176, n27175, n27174, n27173, n27172, 
        n27171, n27170, n27169, n26970;
    wire [31:0]n134;
    
    wire n26969, n26968, n26967, n26966, n26965, n26964, n26963, 
        n26962, n26961, n26960, n26959, n26958, n26957, n26956, 
        n27, n27373, n25, n26, n24, n19, n32, n28, n20, n29, 
        n26_adj_30, n26955;
    
    CCU2D add_19623_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27180), 
          .S0(n7985));
    defparam add_19623_cout.INIT0 = 16'h0000;
    defparam add_19623_cout.INIT1 = 16'h0000;
    defparam add_19623_cout.INJECT1_0 = "NO";
    defparam add_19623_cout.INJECT1_1 = "NO";
    CCU2D add_19623_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27179), .COUT(n27180));
    defparam add_19623_24.INIT0 = 16'h5555;
    defparam add_19623_24.INIT1 = 16'h5555;
    defparam add_19623_24.INJECT1_0 = "NO";
    defparam add_19623_24.INJECT1_1 = "NO";
    CCU2D add_19623_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27178), .COUT(n27179));
    defparam add_19623_22.INIT0 = 16'h5555;
    defparam add_19623_22.INIT1 = 16'h5555;
    defparam add_19623_22.INJECT1_0 = "NO";
    defparam add_19623_22.INJECT1_1 = "NO";
    CCU2D add_19623_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27177), .COUT(n27178));
    defparam add_19623_20.INIT0 = 16'h5555;
    defparam add_19623_20.INIT1 = 16'h5555;
    defparam add_19623_20.INJECT1_0 = "NO";
    defparam add_19623_20.INJECT1_1 = "NO";
    CCU2D add_19623_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27176), .COUT(n27177));
    defparam add_19623_18.INIT0 = 16'h5555;
    defparam add_19623_18.INIT1 = 16'h5555;
    defparam add_19623_18.INJECT1_0 = "NO";
    defparam add_19623_18.INJECT1_1 = "NO";
    CCU2D add_19623_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27175), .COUT(n27176));
    defparam add_19623_16.INIT0 = 16'h5aaa;
    defparam add_19623_16.INIT1 = 16'h5555;
    defparam add_19623_16.INJECT1_0 = "NO";
    defparam add_19623_16.INJECT1_1 = "NO";
    CCU2D add_19623_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27174), .COUT(n27175));
    defparam add_19623_14.INIT0 = 16'h5aaa;
    defparam add_19623_14.INIT1 = 16'h5555;
    defparam add_19623_14.INJECT1_0 = "NO";
    defparam add_19623_14.INJECT1_1 = "NO";
    CCU2D add_19623_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27173), .COUT(n27174));
    defparam add_19623_12.INIT0 = 16'h5555;
    defparam add_19623_12.INIT1 = 16'h5aaa;
    defparam add_19623_12.INJECT1_0 = "NO";
    defparam add_19623_12.INJECT1_1 = "NO";
    CCU2D add_19623_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27172), .COUT(n27173));
    defparam add_19623_10.INIT0 = 16'h5aaa;
    defparam add_19623_10.INIT1 = 16'h5aaa;
    defparam add_19623_10.INJECT1_0 = "NO";
    defparam add_19623_10.INJECT1_1 = "NO";
    CCU2D add_19623_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27171), .COUT(n27172));
    defparam add_19623_8.INIT0 = 16'h5555;
    defparam add_19623_8.INIT1 = 16'h5aaa;
    defparam add_19623_8.INJECT1_0 = "NO";
    defparam add_19623_8.INJECT1_1 = "NO";
    CCU2D add_19623_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27170), .COUT(n27171));
    defparam add_19623_6.INIT0 = 16'h5555;
    defparam add_19623_6.INIT1 = 16'h5555;
    defparam add_19623_6.INJECT1_0 = "NO";
    defparam add_19623_6.INJECT1_1 = "NO";
    CCU2D add_19623_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27169), .COUT(n27170));
    defparam add_19623_4.INIT0 = 16'h5aaa;
    defparam add_19623_4.INIT1 = 16'h5aaa;
    defparam add_19623_4.INJECT1_0 = "NO";
    defparam add_19623_4.INJECT1_1 = "NO";
    CCU2D add_19623_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27169));
    defparam add_19623_2.INIT0 = 16'h7000;
    defparam add_19623_2.INIT1 = 16'h5555;
    defparam add_19623_2.INJECT1_0 = "NO";
    defparam add_19623_2.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26970), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_33.INIT1 = 16'h0000;
    defparam count_2672_add_4_33.INJECT1_0 = "NO";
    defparam count_2672_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26969), .COUT(n26970), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_31.INJECT1_0 = "NO";
    defparam count_2672_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26968), .COUT(n26969), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_29.INJECT1_0 = "NO";
    defparam count_2672_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26967), .COUT(n26968), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_27.INJECT1_0 = "NO";
    defparam count_2672_add_4_27.INJECT1_1 = "NO";
    FD1S3IX clk_o_14 (.D(n7985), .CK(debug_c_c), .CD(n31511), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2672_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26966), .COUT(n26967), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_25.INJECT1_0 = "NO";
    defparam count_2672_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26965), .COUT(n26966), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_23.INJECT1_0 = "NO";
    defparam count_2672_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26964), .COUT(n26965), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_21.INJECT1_0 = "NO";
    defparam count_2672_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26963), .COUT(n26964), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_19.INJECT1_0 = "NO";
    defparam count_2672_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26962), .COUT(n26963), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_17.INJECT1_0 = "NO";
    defparam count_2672_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26961), .COUT(n26962), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_15.INJECT1_0 = "NO";
    defparam count_2672_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26960), .COUT(n26961), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_13.INJECT1_0 = "NO";
    defparam count_2672_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26959), .COUT(n26960), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_11.INJECT1_0 = "NO";
    defparam count_2672_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26958), .COUT(n26959), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_9.INJECT1_0 = "NO";
    defparam count_2672_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26957), .COUT(n26958), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_7.INJECT1_0 = "NO";
    defparam count_2672_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26956), .COUT(n26957), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_5.INJECT1_0 = "NO";
    defparam count_2672_add_4_5.INJECT1_1 = "NO";
    LUT4 i22328_4_lut (.A(n27), .B(n27373), .C(n25), .D(n26), .Z(n29788)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i22328_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n27373)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_30), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_55 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_55.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D count_2672_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26955), .COUT(n26956), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_3.INJECT1_0 = "NO";
    defparam count_2672_add_4_3.INJECT1_1 = "NO";
    LUT4 i12_4_lut_adj_56 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_56.init = 16'h8000;
    CCU2D count_2672_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26955), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672_add_4_1.INIT0 = 16'hF000;
    defparam count_2672_add_4_1.INIT1 = 16'h0555;
    defparam count_2672_add_4_1.INJECT1_0 = "NO";
    defparam count_2672_add_4_1.INJECT1_1 = "NO";
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_30)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    FD1S3IX count_2672__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2875), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i0.GSR = "ENABLED";
    FD1S3IX count_2672__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2875), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i1.GSR = "ENABLED";
    FD1S3IX count_2672__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2875), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i2.GSR = "ENABLED";
    FD1S3IX count_2672__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2875), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i3.GSR = "ENABLED";
    FD1S3IX count_2672__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2875), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i4.GSR = "ENABLED";
    FD1S3IX count_2672__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2875), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i5.GSR = "ENABLED";
    FD1S3IX count_2672__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2875), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i6.GSR = "ENABLED";
    FD1S3IX count_2672__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2875), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i7.GSR = "ENABLED";
    FD1S3IX count_2672__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2875), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i8.GSR = "ENABLED";
    FD1S3IX count_2672__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2875), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i9.GSR = "ENABLED";
    FD1S3IX count_2672__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i10.GSR = "ENABLED";
    FD1S3IX count_2672__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i11.GSR = "ENABLED";
    FD1S3IX count_2672__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i12.GSR = "ENABLED";
    FD1S3IX count_2672__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i13.GSR = "ENABLED";
    FD1S3IX count_2672__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i14.GSR = "ENABLED";
    FD1S3IX count_2672__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i15.GSR = "ENABLED";
    FD1S3IX count_2672__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i16.GSR = "ENABLED";
    FD1S3IX count_2672__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i17.GSR = "ENABLED";
    FD1S3IX count_2672__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i18.GSR = "ENABLED";
    FD1S3IX count_2672__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i19.GSR = "ENABLED";
    FD1S3IX count_2672__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i20.GSR = "ENABLED";
    FD1S3IX count_2672__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i21.GSR = "ENABLED";
    FD1S3IX count_2672__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i22.GSR = "ENABLED";
    FD1S3IX count_2672__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i23.GSR = "ENABLED";
    FD1S3IX count_2672__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i24.GSR = "ENABLED";
    FD1S3IX count_2672__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i25.GSR = "ENABLED";
    FD1S3IX count_2672__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i26.GSR = "ENABLED";
    FD1S3IX count_2672__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i27.GSR = "ENABLED";
    FD1S3IX count_2672__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i28.GSR = "ENABLED";
    FD1S3IX count_2672__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i29.GSR = "ENABLED";
    FD1S3IX count_2672__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i30.GSR = "ENABLED";
    FD1S3IX count_2672__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2875), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2672__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (clk_255kHz, debug_c_c, n241, GND_net, n7916, 
            n31511, n7881, n29831, n14512, n29829, n14513, n2823, 
            n29839, n27540, n29846, n27535, n29817, n13956, n29529, 
            n14, n29943, n14499, n29783, n27563, n29810, n27546, 
            n29826, n27542, n29837, n27549) /* synthesis syn_module_defined=1 */ ;
    output clk_255kHz;
    input debug_c_c;
    input n241;
    input GND_net;
    output n7916;
    input n31511;
    output n7881;
    input n29831;
    output n14512;
    input n29829;
    output n14513;
    input n2823;
    input n29839;
    output n27540;
    input n29846;
    output n27535;
    input n29817;
    output n13956;
    input n29529;
    output n14;
    input n29943;
    output n14499;
    input n29783;
    output n27563;
    input n29810;
    output n27546;
    input n29826;
    output n27542;
    input n29837;
    output n27549;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26714, n26713;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n26712, n26711, n26710, n26709, n26708, n26707, n26706, 
        n26705, n26704, n26703, n26702, n26701, n26700, n26699;
    wire [31:0]n134;
    
    wire n27129, n27128, n27127, n27126, n27125, n27124, n27123, 
        n27122, n27121, n27120, n27119, n27118, n27117, n27116, 
        n27115, n26906, n26905, n26904, n26903, n26902, n26901, 
        n26900, n26899, n26898, n26897, n26896, n26895, n26894, 
        n26893, n26892, n26891;
    
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=538, LSE_RLINE=541 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2058_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26714), .S0(n7916));
    defparam sub_2058_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2058_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2058_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2058_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26713), .COUT(n26714));
    defparam sub_2058_add_2_32.INIT0 = 16'h5555;
    defparam sub_2058_add_2_32.INIT1 = 16'h5555;
    defparam sub_2058_add_2_32.INJECT1_0 = "NO";
    defparam sub_2058_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26712), .COUT(n26713));
    defparam sub_2058_add_2_30.INIT0 = 16'h5555;
    defparam sub_2058_add_2_30.INIT1 = 16'h5555;
    defparam sub_2058_add_2_30.INJECT1_0 = "NO";
    defparam sub_2058_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26711), .COUT(n26712));
    defparam sub_2058_add_2_28.INIT0 = 16'h5555;
    defparam sub_2058_add_2_28.INIT1 = 16'h5555;
    defparam sub_2058_add_2_28.INJECT1_0 = "NO";
    defparam sub_2058_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26710), .COUT(n26711));
    defparam sub_2058_add_2_26.INIT0 = 16'h5555;
    defparam sub_2058_add_2_26.INIT1 = 16'h5555;
    defparam sub_2058_add_2_26.INJECT1_0 = "NO";
    defparam sub_2058_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26709), .COUT(n26710));
    defparam sub_2058_add_2_24.INIT0 = 16'h5555;
    defparam sub_2058_add_2_24.INIT1 = 16'h5555;
    defparam sub_2058_add_2_24.INJECT1_0 = "NO";
    defparam sub_2058_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26708), .COUT(n26709));
    defparam sub_2058_add_2_22.INIT0 = 16'h5555;
    defparam sub_2058_add_2_22.INIT1 = 16'h5555;
    defparam sub_2058_add_2_22.INJECT1_0 = "NO";
    defparam sub_2058_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26707), .COUT(n26708));
    defparam sub_2058_add_2_20.INIT0 = 16'h5555;
    defparam sub_2058_add_2_20.INIT1 = 16'h5555;
    defparam sub_2058_add_2_20.INJECT1_0 = "NO";
    defparam sub_2058_add_2_20.INJECT1_1 = "NO";
    LUT4 i22372_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29831), 
         .Z(n14512)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22372_2_lut_4_lut.init = 16'h1000;
    LUT4 i22370_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29829), 
         .Z(n14513)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22370_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_2058_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26706), .COUT(n26707));
    defparam sub_2058_add_2_18.INIT0 = 16'h5555;
    defparam sub_2058_add_2_18.INIT1 = 16'h5555;
    defparam sub_2058_add_2_18.INJECT1_0 = "NO";
    defparam sub_2058_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26705), .COUT(n26706));
    defparam sub_2058_add_2_16.INIT0 = 16'h5555;
    defparam sub_2058_add_2_16.INIT1 = 16'h5555;
    defparam sub_2058_add_2_16.INJECT1_0 = "NO";
    defparam sub_2058_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26704), .COUT(n26705));
    defparam sub_2058_add_2_14.INIT0 = 16'h5555;
    defparam sub_2058_add_2_14.INIT1 = 16'h5555;
    defparam sub_2058_add_2_14.INJECT1_0 = "NO";
    defparam sub_2058_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26703), .COUT(n26704));
    defparam sub_2058_add_2_12.INIT0 = 16'h5555;
    defparam sub_2058_add_2_12.INIT1 = 16'h5555;
    defparam sub_2058_add_2_12.INJECT1_0 = "NO";
    defparam sub_2058_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26702), .COUT(n26703));
    defparam sub_2058_add_2_10.INIT0 = 16'h5555;
    defparam sub_2058_add_2_10.INIT1 = 16'h5555;
    defparam sub_2058_add_2_10.INJECT1_0 = "NO";
    defparam sub_2058_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26701), .COUT(n26702));
    defparam sub_2058_add_2_8.INIT0 = 16'h5555;
    defparam sub_2058_add_2_8.INIT1 = 16'h5555;
    defparam sub_2058_add_2_8.INJECT1_0 = "NO";
    defparam sub_2058_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26700), .COUT(n26701));
    defparam sub_2058_add_2_6.INIT0 = 16'h5555;
    defparam sub_2058_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_2058_add_2_6.INJECT1_0 = "NO";
    defparam sub_2058_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2058_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26699), .COUT(n26700));
    defparam sub_2058_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2058_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_2058_add_2_4.INJECT1_0 = "NO";
    defparam sub_2058_add_2_4.INJECT1_1 = "NO";
    FD1S3IX count_2670__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2823), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i0.GSR = "ENABLED";
    CCU2D sub_2058_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26699));
    defparam sub_2058_add_2_2.INIT0 = 16'h0000;
    defparam sub_2058_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2058_add_2_2.INJECT1_0 = "NO";
    defparam sub_2058_add_2_2.INJECT1_1 = "NO";
    LUT4 i22380_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29839), 
         .Z(n27540)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22380_2_lut_4_lut.init = 16'h1000;
    CCU2D add_19626_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27129), 
          .S1(n7881));
    defparam add_19626_32.INIT0 = 16'h5555;
    defparam add_19626_32.INIT1 = 16'h0000;
    defparam add_19626_32.INJECT1_0 = "NO";
    defparam add_19626_32.INJECT1_1 = "NO";
    CCU2D add_19626_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27128), .COUT(n27129));
    defparam add_19626_30.INIT0 = 16'h5555;
    defparam add_19626_30.INIT1 = 16'h5555;
    defparam add_19626_30.INJECT1_0 = "NO";
    defparam add_19626_30.INJECT1_1 = "NO";
    CCU2D add_19626_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27127), .COUT(n27128));
    defparam add_19626_28.INIT0 = 16'h5555;
    defparam add_19626_28.INIT1 = 16'h5555;
    defparam add_19626_28.INJECT1_0 = "NO";
    defparam add_19626_28.INJECT1_1 = "NO";
    CCU2D add_19626_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27126), .COUT(n27127));
    defparam add_19626_26.INIT0 = 16'h5555;
    defparam add_19626_26.INIT1 = 16'h5555;
    defparam add_19626_26.INJECT1_0 = "NO";
    defparam add_19626_26.INJECT1_1 = "NO";
    LUT4 i22387_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29846), 
         .Z(n27535)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22387_2_lut_4_lut.init = 16'h1000;
    CCU2D add_19626_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27125), .COUT(n27126));
    defparam add_19626_24.INIT0 = 16'h5555;
    defparam add_19626_24.INIT1 = 16'h5555;
    defparam add_19626_24.INJECT1_0 = "NO";
    defparam add_19626_24.INJECT1_1 = "NO";
    LUT4 i22358_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29817), 
         .Z(n13956)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22358_2_lut_4_lut.init = 16'h1000;
    LUT4 i5_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29529), 
         .Z(n14)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i5_2_lut_4_lut.init = 16'h0010;
    LUT4 i22484_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29943), 
         .Z(n14499)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22484_2_lut_4_lut.init = 16'h1000;
    CCU2D add_19626_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27124), .COUT(n27125));
    defparam add_19626_22.INIT0 = 16'h5555;
    defparam add_19626_22.INIT1 = 16'h5555;
    defparam add_19626_22.INJECT1_0 = "NO";
    defparam add_19626_22.INJECT1_1 = "NO";
    CCU2D add_19626_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27123), .COUT(n27124));
    defparam add_19626_20.INIT0 = 16'h5555;
    defparam add_19626_20.INIT1 = 16'h5555;
    defparam add_19626_20.INJECT1_0 = "NO";
    defparam add_19626_20.INJECT1_1 = "NO";
    CCU2D add_19626_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27122), .COUT(n27123));
    defparam add_19626_18.INIT0 = 16'h5555;
    defparam add_19626_18.INIT1 = 16'h5555;
    defparam add_19626_18.INJECT1_0 = "NO";
    defparam add_19626_18.INJECT1_1 = "NO";
    CCU2D add_19626_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27121), .COUT(n27122));
    defparam add_19626_16.INIT0 = 16'h5555;
    defparam add_19626_16.INIT1 = 16'h5555;
    defparam add_19626_16.INJECT1_0 = "NO";
    defparam add_19626_16.INJECT1_1 = "NO";
    CCU2D add_19626_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27120), .COUT(n27121));
    defparam add_19626_14.INIT0 = 16'h5555;
    defparam add_19626_14.INIT1 = 16'h5555;
    defparam add_19626_14.INJECT1_0 = "NO";
    defparam add_19626_14.INJECT1_1 = "NO";
    CCU2D add_19626_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27119), .COUT(n27120));
    defparam add_19626_12.INIT0 = 16'h5555;
    defparam add_19626_12.INIT1 = 16'h5555;
    defparam add_19626_12.INJECT1_0 = "NO";
    defparam add_19626_12.INJECT1_1 = "NO";
    CCU2D add_19626_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27118), .COUT(n27119));
    defparam add_19626_10.INIT0 = 16'h5555;
    defparam add_19626_10.INIT1 = 16'h5555;
    defparam add_19626_10.INJECT1_0 = "NO";
    defparam add_19626_10.INJECT1_1 = "NO";
    CCU2D add_19626_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27117), 
          .COUT(n27118));
    defparam add_19626_8.INIT0 = 16'h5555;
    defparam add_19626_8.INIT1 = 16'h5555;
    defparam add_19626_8.INJECT1_0 = "NO";
    defparam add_19626_8.INJECT1_1 = "NO";
    CCU2D add_19626_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27116), 
          .COUT(n27117));
    defparam add_19626_6.INIT0 = 16'h5555;
    defparam add_19626_6.INIT1 = 16'h5555;
    defparam add_19626_6.INJECT1_0 = "NO";
    defparam add_19626_6.INJECT1_1 = "NO";
    CCU2D add_19626_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27115), 
          .COUT(n27116));
    defparam add_19626_4.INIT0 = 16'h5555;
    defparam add_19626_4.INIT1 = 16'h5aaa;
    defparam add_19626_4.INJECT1_0 = "NO";
    defparam add_19626_4.INJECT1_1 = "NO";
    CCU2D add_19626_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27115));
    defparam add_19626_2.INIT0 = 16'h7000;
    defparam add_19626_2.INIT1 = 16'h5aaa;
    defparam add_19626_2.INJECT1_0 = "NO";
    defparam add_19626_2.INJECT1_1 = "NO";
    LUT4 i22324_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29783), 
         .Z(n27563)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22324_2_lut_4_lut.init = 16'h1000;
    LUT4 i22351_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29810), 
         .Z(n27546)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22351_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2670_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26906), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_33.INIT1 = 16'h0000;
    defparam count_2670_add_4_33.INJECT1_0 = "NO";
    defparam count_2670_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26905), .COUT(n26906), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_31.INJECT1_0 = "NO";
    defparam count_2670_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26904), .COUT(n26905), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_29.INJECT1_0 = "NO";
    defparam count_2670_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26903), .COUT(n26904), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_27.INJECT1_0 = "NO";
    defparam count_2670_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26902), .COUT(n26903), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_25.INJECT1_0 = "NO";
    defparam count_2670_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26901), .COUT(n26902), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_23.INJECT1_0 = "NO";
    defparam count_2670_add_4_23.INJECT1_1 = "NO";
    FD1S3IX count_2670__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2823), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i1.GSR = "ENABLED";
    FD1S3IX count_2670__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2823), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i2.GSR = "ENABLED";
    FD1S3IX count_2670__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2823), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i3.GSR = "ENABLED";
    FD1S3IX count_2670__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2823), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i4.GSR = "ENABLED";
    FD1S3IX count_2670__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2823), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i5.GSR = "ENABLED";
    FD1S3IX count_2670__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2823), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i6.GSR = "ENABLED";
    FD1S3IX count_2670__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2823), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i7.GSR = "ENABLED";
    FD1S3IX count_2670__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2823), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i8.GSR = "ENABLED";
    FD1S3IX count_2670__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2823), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i9.GSR = "ENABLED";
    FD1S3IX count_2670__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i10.GSR = "ENABLED";
    FD1S3IX count_2670__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i11.GSR = "ENABLED";
    FD1S3IX count_2670__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i12.GSR = "ENABLED";
    FD1S3IX count_2670__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i13.GSR = "ENABLED";
    FD1S3IX count_2670__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i14.GSR = "ENABLED";
    FD1S3IX count_2670__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i15.GSR = "ENABLED";
    FD1S3IX count_2670__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i16.GSR = "ENABLED";
    FD1S3IX count_2670__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i17.GSR = "ENABLED";
    FD1S3IX count_2670__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i18.GSR = "ENABLED";
    FD1S3IX count_2670__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i19.GSR = "ENABLED";
    FD1S3IX count_2670__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i20.GSR = "ENABLED";
    FD1S3IX count_2670__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i21.GSR = "ENABLED";
    FD1S3IX count_2670__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i22.GSR = "ENABLED";
    FD1S3IX count_2670__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i23.GSR = "ENABLED";
    FD1S3IX count_2670__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i24.GSR = "ENABLED";
    FD1S3IX count_2670__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i25.GSR = "ENABLED";
    FD1S3IX count_2670__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i26.GSR = "ENABLED";
    FD1S3IX count_2670__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i27.GSR = "ENABLED";
    FD1S3IX count_2670__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i28.GSR = "ENABLED";
    FD1S3IX count_2670__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i29.GSR = "ENABLED";
    FD1S3IX count_2670__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i30.GSR = "ENABLED";
    FD1S3IX count_2670__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2823), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670__i31.GSR = "ENABLED";
    CCU2D count_2670_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26900), .COUT(n26901), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_21.INJECT1_0 = "NO";
    defparam count_2670_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26899), .COUT(n26900), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_19.INJECT1_0 = "NO";
    defparam count_2670_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26898), .COUT(n26899), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_17.INJECT1_0 = "NO";
    defparam count_2670_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26897), .COUT(n26898), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_15.INJECT1_0 = "NO";
    defparam count_2670_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26896), .COUT(n26897), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_13.INJECT1_0 = "NO";
    defparam count_2670_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26895), .COUT(n26896), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_11.INJECT1_0 = "NO";
    defparam count_2670_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26894), .COUT(n26895), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_9.INJECT1_0 = "NO";
    defparam count_2670_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26893), .COUT(n26894), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_7.INJECT1_0 = "NO";
    defparam count_2670_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26892), .COUT(n26893), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_5.INJECT1_0 = "NO";
    defparam count_2670_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26891), .COUT(n26892), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2670_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2670_add_4_3.INJECT1_0 = "NO";
    defparam count_2670_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2670_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26891), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2670_add_4_1.INIT0 = 16'hF000;
    defparam count_2670_add_4_1.INIT1 = 16'h0555;
    defparam count_2670_add_4_1.INJECT1_0 = "NO";
    defparam count_2670_add_4_1.INJECT1_1 = "NO";
    LUT4 i22367_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29826), 
         .Z(n27542)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22367_2_lut_4_lut.init = 16'h1000;
    LUT4 i22378_2_lut_4_lut (.A(n31511), .B(clk_255kHz), .C(n7881), .D(n29837), 
         .Z(n27549)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22378_2_lut_4_lut.init = 16'h1000;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (debug_c_c, n31511, databus, n4180, 
            \read_size[0] , n13940, n9378, Stepper_X_M0_c_0, n13916, 
            prev_step_clk, step_clk, limit_latched, prev_limit_latched, 
            n9296, prev_select, n31473, \register_addr[1] , Stepper_X_Dir_c, 
            \register_addr[0] , n1, Stepper_X_En_c, Stepper_X_M1_c_1, 
            \control_reg[7] , n12158, Stepper_X_M2_c_2, \read_size[2] , 
            n31434, n34, n27444, n29136, limit_c_0, read_value, 
            n31424, n24, n31420, VCC_net, GND_net, Stepper_X_nFault_c, 
            Stepper_X_Step_c, n31408, n8055, n8089, n17034) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31511;
    input [31:0]databus;
    input n4180;
    output \read_size[0] ;
    input n13940;
    input n9378;
    output Stepper_X_M0_c_0;
    input n13916;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    input n9296;
    output prev_select;
    input n31473;
    input \register_addr[1] ;
    output Stepper_X_Dir_c;
    input \register_addr[0] ;
    input n1;
    output Stepper_X_En_c;
    output Stepper_X_M1_c_1;
    output \control_reg[7] ;
    input n12158;
    output Stepper_X_M2_c_2;
    output \read_size[2] ;
    input n31434;
    input n34;
    output n27444;
    input n29136;
    input limit_c_0;
    output [31:0]read_value;
    input n31424;
    input n24;
    input n31420;
    input VCC_net;
    input GND_net;
    input Stepper_X_nFault_c;
    output Stepper_X_Step_c;
    input n31408;
    output n8055;
    output n8089;
    input n17034;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n4181;
    wire [31:0]n224;
    
    wire n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n1_c, n2;
    wire [31:0]n6498;
    
    wire n29695, n29696, n1_adj_22, n2_adj_23, n2_adj_25;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n1_adj_26, n29683, n29684, n29685, n2_adj_27, fault_latched, 
        n29764, n29765, n49, n62, n58, n50, n41, n60, n54, 
        n42, n52, n38, n56, n46, n29697, n1_adj_28, n2_adj_29, 
        n29766, n29141, n29143, n29144, n29146, n29142, n29147, 
        n29148, n29150, n29145, n29151, n29149, n29152, n29153, 
        n29154, n29155, n29139, n29137, n29140, n29157, n29158, 
        n29159, n29160, n29138, n29156, int_step, n26882, n26881, 
        n26880, n26879, n26878, n26877, n26876, n26875, n26874, 
        n26873, n26872, n26871, n26870, n26869, n26868, n26867;
    
    FD1S3IX steps_reg__i26 (.D(n4181[26]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4181[25]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4181[24]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4181[23]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4181[22]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4181[21]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4181[20]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4181[19]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4181[18]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4181[17]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4181[16]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4181[15]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4181[14]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4181[13]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4181[12]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4181[11]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4181[10]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4181[9]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4181[8]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4181[7]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4181[6]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4181[5]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4181[4]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4181[3]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4181[2]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4181[1]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1621_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4180), .Z(n4181[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i10_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i0 (.D(n4181[0]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n9378), .SP(n13940), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n13916), .CD(n31511), 
            .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31473), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 mux_1621_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4180), .Z(n4181[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i9_3_lut.init = 16'hcaca;
    PFUMX mux_1929_Mux_5_i3 (.BLUT(n1_c), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n6498[5]));
    LUT4 i22135_3_lut (.A(Stepper_X_M0_c_0), .B(div_factor_reg[0]), .C(\register_addr[1] ), 
         .Z(n29695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22135_3_lut.init = 16'hcaca;
    LUT4 i22136_3_lut (.A(limit_latched), .B(steps_reg[0]), .C(\register_addr[1] ), 
         .Z(n29696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22136_3_lut.init = 16'hcaca;
    LUT4 i15138_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_c)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15138_2_lut.init = 16'h2222;
    LUT4 mux_1929_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1929_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4180), .Z(n4181[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i8_3_lut.init = 16'hcaca;
    PFUMX mux_1929_Mux_6_i3 (.BLUT(n1_adj_22), .ALUT(n2_adj_23), .C0(\register_addr[1] ), 
          .Z(n6498[6]));
    LUT4 mux_1621_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4180), .Z(n4181[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i7_3_lut.init = 16'hcaca;
    PFUMX mux_1929_Mux_7_i3 (.BLUT(n1), .ALUT(n2_adj_25), .C0(\register_addr[1] ), 
          .Z(n6498[7]));
    LUT4 mux_1621_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4180), 
         .Z(n4181[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4180), .Z(n4181[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4180), .Z(n4181[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4180), 
         .Z(n4181[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4180), 
         .Z(n4181[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4180), .Z(n4181[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4180), 
         .Z(n4181[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4180), .Z(n4181[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4180), .Z(n4181[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4180), 
         .Z(n4181[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4180), 
         .Z(n4181[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4180), 
         .Z(n4181[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4180), 
         .Z(n4181[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i13_3_lut.init = 16'hcaca;
    LUT4 i15135_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_22)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15135_2_lut.init = 16'h2222;
    LUT4 mux_1929_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1929_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1929_Mux_7_i2_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), 
         .C(\register_addr[0] ), .Z(n2_adj_25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1929_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4180), 
         .Z(n4181[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4180), 
         .Z(n4181[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i11_3_lut.init = 16'hcaca;
    LUT4 i15140_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1_adj_26)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15140_2_lut.init = 16'h2222;
    PFUMX i22125 (.BLUT(n29683), .ALUT(n29684), .C0(\register_addr[1] ), 
          .Z(n29685));
    LUT4 mux_1929_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2_adj_27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1929_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i22204_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22204_3_lut.init = 16'hcaca;
    LUT4 i22205_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22205_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4180), 
         .Z(n4181[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4180), 
         .Z(n4181[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i17_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9296), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9296), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9296), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9296), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9296), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9296), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9296), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n9296), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13916), .CD(n12158), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13916), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13916), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13916), .CD(n31511), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13916), .PD(n31511), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13916), .CD(n31511), 
            .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13916), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n31434), .SP(n13940), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 mux_1621_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4180), 
         .Z(n4181[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i21_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i31 (.D(n4181[31]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4181[30]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4181[29]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4181[28]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    LUT4 i22123_3_lut (.A(Stepper_X_M2_c_2), .B(n34), .C(\register_addr[0] ), 
         .Z(n29683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22123_3_lut.init = 16'hcaca;
    LUT4 i22124_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n29684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22124_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27444)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 mux_1621_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4180), 
         .Z(n4181[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4180), 
         .Z(n4181[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4180), 
         .Z(n4181[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i29_3_lut.init = 16'hcaca;
    LUT4 i17_4_lut (.A(steps_reg[8]), .B(steps_reg[27]), .C(steps_reg[31]), 
         .D(steps_reg[30]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[15]), .B(n52), .C(n38), .D(steps_reg[11]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[20]), .B(steps_reg[18]), .C(steps_reg[24]), 
         .D(steps_reg[4]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[9]), .B(steps_reg[12]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[5]), .B(n56), .C(n46), .D(steps_reg[6]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[7]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[16]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[17]), .B(steps_reg[21]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    PFUMX i22137 (.BLUT(n29695), .ALUT(n29696), .C0(\register_addr[0] ), 
          .Z(n29697));
    LUT4 mux_1621_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4180), 
         .Z(n4181[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i15_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i27 (.D(n4181[27]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    LUT4 i24_4_lut (.A(steps_reg[19]), .B(steps_reg[3]), .C(steps_reg[22]), 
         .D(steps_reg[13]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[10]), .B(steps_reg[14]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[29]), .B(steps_reg[0]), .C(steps_reg[2]), 
         .D(steps_reg[1]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[28]), .B(steps_reg[23]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1621_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4180), .Z(n4181[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i1_3_lut.init = 16'hcaca;
    LUT4 i15139_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_28)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15139_2_lut.init = 16'h2222;
    LUT4 mux_1929_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2_adj_29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1929_Mux_4_i2_3_lut.init = 16'hcaca;
    PFUMX mux_1929_Mux_3_i3 (.BLUT(n1_adj_26), .ALUT(n2_adj_27), .C0(\register_addr[1] ), 
          .Z(n6498[3]));
    PFUMX i22206 (.BLUT(n29764), .ALUT(n29765), .C0(\register_addr[1] ), 
          .Z(n29766));
    LUT4 i1_4_lut (.A(div_factor_reg[31]), .B(n29136), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n29141)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hc088;
    LUT4 mux_1621_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4180), 
         .Z(n4181[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i20_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_32 (.A(div_factor_reg[30]), .B(n29136), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29143)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_32.init = 16'hc088;
    LUT4 i1_4_lut_adj_33 (.A(div_factor_reg[29]), .B(n29136), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29144)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_33.init = 16'hc088;
    LUT4 i1_4_lut_adj_34 (.A(div_factor_reg[28]), .B(n29136), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n29146)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_34.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_35 (.A(div_factor_reg[27]), .B(n29136), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n29142)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_35.init = 16'hc088;
    FD1P3AX read_value__i31 (.D(n29141), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29143), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29144), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29146), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29142), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29147), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29148), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29150), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29145), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29151), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29149), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29152), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    LUT4 mux_1621_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4180), 
         .Z(n4181[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i16_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i19 (.D(n29153), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29154), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29155), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29139), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29137), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29140), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29157), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29158), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29159), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29160), .SP(n13940), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29138), .SP(n13940), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29156), .SP(n13940), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6498[7]), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6498[6]), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6498[5]), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6498[4]), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6498[3]), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29685), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29766), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_36 (.A(div_factor_reg[26]), .B(n29136), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n29147)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_36.init = 16'hc088;
    FD1P3AX int_step_182 (.D(n31420), .SP(n24), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_37 (.A(div_factor_reg[25]), .B(n29136), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n29148)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_37.init = 16'hc088;
    LUT4 i1_4_lut_adj_38 (.A(div_factor_reg[24]), .B(n29136), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n29150)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_38.init = 16'hc088;
    LUT4 i1_4_lut_adj_39 (.A(div_factor_reg[23]), .B(n29136), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n29145)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_39.init = 16'hc088;
    LUT4 i1_4_lut_adj_40 (.A(div_factor_reg[22]), .B(n29136), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n29151)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_40.init = 16'hc088;
    LUT4 i1_4_lut_adj_41 (.A(div_factor_reg[21]), .B(n29136), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n29149)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_41.init = 16'hc088;
    LUT4 i1_4_lut_adj_42 (.A(div_factor_reg[20]), .B(n29136), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n29152)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_42.init = 16'hc088;
    LUT4 i1_4_lut_adj_43 (.A(div_factor_reg[19]), .B(n29136), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n29153)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_43.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26882), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_44 (.A(div_factor_reg[18]), .B(n29136), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n29154)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_44.init = 16'hc088;
    LUT4 i1_4_lut_adj_45 (.A(div_factor_reg[17]), .B(n29136), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n29155)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_45.init = 16'hc088;
    LUT4 i1_4_lut_adj_46 (.A(div_factor_reg[16]), .B(n29136), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n29139)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_46.init = 16'hc088;
    LUT4 i1_4_lut_adj_47 (.A(div_factor_reg[15]), .B(n29136), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n29137)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_47.init = 16'hc088;
    LUT4 i1_4_lut_adj_48 (.A(div_factor_reg[14]), .B(n29136), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n29140)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_48.init = 16'hc088;
    LUT4 i1_4_lut_adj_49 (.A(div_factor_reg[13]), .B(n29136), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n29157)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_49.init = 16'hc088;
    LUT4 i1_4_lut_adj_50 (.A(div_factor_reg[12]), .B(n29136), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n29158)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_50.init = 16'hc088;
    LUT4 i1_4_lut_adj_51 (.A(div_factor_reg[11]), .B(n29136), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n29159)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_51.init = 16'hc088;
    LUT4 i1_4_lut_adj_52 (.A(div_factor_reg[10]), .B(n29136), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n29160)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_52.init = 16'hc088;
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26881), .COUT(n26882), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_53 (.A(div_factor_reg[9]), .B(n29136), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n29138)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_53.init = 16'hc088;
    LUT4 i1_4_lut_adj_54 (.A(div_factor_reg[8]), .B(n29136), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29156)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_54.init = 16'hc088;
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26880), .COUT(n26881), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26879), .COUT(n26880), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26878), .COUT(n26879), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26877), .COUT(n26878), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    FD1P3IX read_value__i0 (.D(n29697), .SP(n13940), .CD(n31424), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=578, LSE_RLINE=591 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26876), .COUT(n26877), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26875), .COUT(n26876), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26874), .COUT(n26875), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26873), .COUT(n26874), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26872), .COUT(n26873), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26871), .COUT(n26872), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26870), .COUT(n26871), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26869), .COUT(n26870), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26868), .COUT(n26869), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 mux_1621_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4180), 
         .Z(n4181[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i19_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26867), .COUT(n26868), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n34), .D1(prev_step_clk), 
          .COUT(n26867), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    PFUMX mux_1929_Mux_4_i3 (.BLUT(n1_adj_28), .ALUT(n2_adj_29), .C0(\register_addr[1] ), 
          .Z(n6498[4]));
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1621_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4180), 
         .Z(n4181[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1621_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4180), 
         .Z(n4181[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1621_i25_3_lut.init = 16'hcaca;
    ClockDivider_U8 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n31511(n31511), .n31408(n31408), .n8055(n8055), 
            .div_factor_reg({div_factor_reg}), .n8089(n8089), .n17034(n17034)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (GND_net, step_clk, debug_c_c, n31511, n31408, 
            n8055, div_factor_reg, n8089, n17034) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31511;
    input n31408;
    output n8055;
    input [31:0]div_factor_reg;
    output n8089;
    input n17034;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26995;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n26996, n26994, n26993, n26992, n26991, n26990, n26989, 
        n26988, n26987, n8020, n26818;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n26817, n26698, n26816, n26697, n26696, n26695, n26815, 
        n26814, n26813, n26812, n26811, n26810, n26694, n26693, 
        n26809, n26808, n26692, n26807, n26806, n26805, n26691, 
        n26804, n26690, n26803, n26689, n26688, n26687, n26686, 
        n26685, n26684, n26683, n26682, n26681, n26680, n26679, 
        n26678, n26677, n26676, n26675, n26674, n26673, n26672, 
        n26671, n26670, n26669, n26668, n26667, n26666, n26665, 
        n26664, n26663, n26662, n26661, n26660, n26659, n26658, 
        n26657, n26656, n26655, n26654, n26653, n26652, n26651, 
        n27002, n27001, n27000, n26999, n26998, n26997;
    
    CCU2D count_2673_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26995), .COUT(n26996), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_19.INJECT1_0 = "NO";
    defparam count_2673_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26994), .COUT(n26995), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_17.INJECT1_0 = "NO";
    defparam count_2673_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26993), .COUT(n26994), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_15.INJECT1_0 = "NO";
    defparam count_2673_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26992), .COUT(n26993), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_13.INJECT1_0 = "NO";
    defparam count_2673_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26991), .COUT(n26992), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_11.INJECT1_0 = "NO";
    defparam count_2673_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26990), .COUT(n26991), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_9.INJECT1_0 = "NO";
    defparam count_2673_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26989), .COUT(n26990), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_7.INJECT1_0 = "NO";
    defparam count_2673_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26988), .COUT(n26989), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_5.INJECT1_0 = "NO";
    defparam count_2673_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26987), .COUT(n26988), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_3.INJECT1_0 = "NO";
    defparam count_2673_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26987), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_1.INIT0 = 16'hF000;
    defparam count_2673_add_4_1.INIT1 = 16'h0555;
    defparam count_2673_add_4_1.INJECT1_0 = "NO";
    defparam count_2673_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8020), .CK(debug_c_c), .CD(n31511), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26818), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26817), .COUT(n26818), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26698), .S1(n8020));
    defparam sub_2063_add_2_33.INIT0 = 16'h5555;
    defparam sub_2063_add_2_33.INIT1 = 16'h0000;
    defparam sub_2063_add_2_33.INJECT1_0 = "NO";
    defparam sub_2063_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26816), .COUT(n26817), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26697), .COUT(n26698));
    defparam sub_2063_add_2_31.INIT0 = 16'h5999;
    defparam sub_2063_add_2_31.INIT1 = 16'h5999;
    defparam sub_2063_add_2_31.INJECT1_0 = "NO";
    defparam sub_2063_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26696), .COUT(n26697));
    defparam sub_2063_add_2_29.INIT0 = 16'h5999;
    defparam sub_2063_add_2_29.INIT1 = 16'h5999;
    defparam sub_2063_add_2_29.INJECT1_0 = "NO";
    defparam sub_2063_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26695), .COUT(n26696));
    defparam sub_2063_add_2_27.INIT0 = 16'h5999;
    defparam sub_2063_add_2_27.INIT1 = 16'h5999;
    defparam sub_2063_add_2_27.INJECT1_0 = "NO";
    defparam sub_2063_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26815), .COUT(n26816), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26814), .COUT(n26815), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26813), .COUT(n26814), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26812), .COUT(n26813), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26811), .COUT(n26812), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26810), .COUT(n26811), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26694), .COUT(n26695));
    defparam sub_2063_add_2_25.INIT0 = 16'h5999;
    defparam sub_2063_add_2_25.INIT1 = 16'h5999;
    defparam sub_2063_add_2_25.INJECT1_0 = "NO";
    defparam sub_2063_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26693), .COUT(n26694));
    defparam sub_2063_add_2_23.INIT0 = 16'h5999;
    defparam sub_2063_add_2_23.INIT1 = 16'h5999;
    defparam sub_2063_add_2_23.INJECT1_0 = "NO";
    defparam sub_2063_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26809), .COUT(n26810), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26808), .COUT(n26809), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26692), .COUT(n26693));
    defparam sub_2063_add_2_21.INIT0 = 16'h5999;
    defparam sub_2063_add_2_21.INIT1 = 16'h5999;
    defparam sub_2063_add_2_21.INJECT1_0 = "NO";
    defparam sub_2063_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26807), .COUT(n26808), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26806), .COUT(n26807), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26805), .COUT(n26806), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26691), .COUT(n26692));
    defparam sub_2063_add_2_19.INIT0 = 16'h5999;
    defparam sub_2063_add_2_19.INIT1 = 16'h5999;
    defparam sub_2063_add_2_19.INJECT1_0 = "NO";
    defparam sub_2063_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26804), .COUT(n26805), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26690), .COUT(n26691));
    defparam sub_2063_add_2_17.INIT0 = 16'h5999;
    defparam sub_2063_add_2_17.INIT1 = 16'h5999;
    defparam sub_2063_add_2_17.INJECT1_0 = "NO";
    defparam sub_2063_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26803), .COUT(n26804), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26803), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26689), .COUT(n26690));
    defparam sub_2063_add_2_15.INIT0 = 16'h5999;
    defparam sub_2063_add_2_15.INIT1 = 16'h5999;
    defparam sub_2063_add_2_15.INJECT1_0 = "NO";
    defparam sub_2063_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26688), .COUT(n26689));
    defparam sub_2063_add_2_13.INIT0 = 16'h5999;
    defparam sub_2063_add_2_13.INIT1 = 16'h5999;
    defparam sub_2063_add_2_13.INJECT1_0 = "NO";
    defparam sub_2063_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26687), .COUT(n26688));
    defparam sub_2063_add_2_11.INIT0 = 16'h5999;
    defparam sub_2063_add_2_11.INIT1 = 16'h5999;
    defparam sub_2063_add_2_11.INJECT1_0 = "NO";
    defparam sub_2063_add_2_11.INJECT1_1 = "NO";
    FD1S3IX count_2673__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i0.GSR = "ENABLED";
    CCU2D sub_2063_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26686), .COUT(n26687));
    defparam sub_2063_add_2_9.INIT0 = 16'h5999;
    defparam sub_2063_add_2_9.INIT1 = 16'h5999;
    defparam sub_2063_add_2_9.INJECT1_0 = "NO";
    defparam sub_2063_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26685), .COUT(n26686));
    defparam sub_2063_add_2_7.INIT0 = 16'h5999;
    defparam sub_2063_add_2_7.INIT1 = 16'h5999;
    defparam sub_2063_add_2_7.INJECT1_0 = "NO";
    defparam sub_2063_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26684), .COUT(n26685));
    defparam sub_2063_add_2_5.INIT0 = 16'h5999;
    defparam sub_2063_add_2_5.INIT1 = 16'h5999;
    defparam sub_2063_add_2_5.INJECT1_0 = "NO";
    defparam sub_2063_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26683), .COUT(n26684));
    defparam sub_2063_add_2_3.INIT0 = 16'h5999;
    defparam sub_2063_add_2_3.INIT1 = 16'h5999;
    defparam sub_2063_add_2_3.INJECT1_0 = "NO";
    defparam sub_2063_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2063_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26683));
    defparam sub_2063_add_2_1.INIT0 = 16'h0000;
    defparam sub_2063_add_2_1.INIT1 = 16'h5999;
    defparam sub_2063_add_2_1.INJECT1_0 = "NO";
    defparam sub_2063_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26682), .S1(n8055));
    defparam sub_2065_add_2_33.INIT0 = 16'h5999;
    defparam sub_2065_add_2_33.INIT1 = 16'h0000;
    defparam sub_2065_add_2_33.INJECT1_0 = "NO";
    defparam sub_2065_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26681), .COUT(n26682));
    defparam sub_2065_add_2_31.INIT0 = 16'h5999;
    defparam sub_2065_add_2_31.INIT1 = 16'h5999;
    defparam sub_2065_add_2_31.INJECT1_0 = "NO";
    defparam sub_2065_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26680), .COUT(n26681));
    defparam sub_2065_add_2_29.INIT0 = 16'h5999;
    defparam sub_2065_add_2_29.INIT1 = 16'h5999;
    defparam sub_2065_add_2_29.INJECT1_0 = "NO";
    defparam sub_2065_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26679), .COUT(n26680));
    defparam sub_2065_add_2_27.INIT0 = 16'h5999;
    defparam sub_2065_add_2_27.INIT1 = 16'h5999;
    defparam sub_2065_add_2_27.INJECT1_0 = "NO";
    defparam sub_2065_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26678), .COUT(n26679));
    defparam sub_2065_add_2_25.INIT0 = 16'h5999;
    defparam sub_2065_add_2_25.INIT1 = 16'h5999;
    defparam sub_2065_add_2_25.INJECT1_0 = "NO";
    defparam sub_2065_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26677), .COUT(n26678));
    defparam sub_2065_add_2_23.INIT0 = 16'h5999;
    defparam sub_2065_add_2_23.INIT1 = 16'h5999;
    defparam sub_2065_add_2_23.INJECT1_0 = "NO";
    defparam sub_2065_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26676), .COUT(n26677));
    defparam sub_2065_add_2_21.INIT0 = 16'h5999;
    defparam sub_2065_add_2_21.INIT1 = 16'h5999;
    defparam sub_2065_add_2_21.INJECT1_0 = "NO";
    defparam sub_2065_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26675), .COUT(n26676));
    defparam sub_2065_add_2_19.INIT0 = 16'h5999;
    defparam sub_2065_add_2_19.INIT1 = 16'h5999;
    defparam sub_2065_add_2_19.INJECT1_0 = "NO";
    defparam sub_2065_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26674), .COUT(n26675));
    defparam sub_2065_add_2_17.INIT0 = 16'h5999;
    defparam sub_2065_add_2_17.INIT1 = 16'h5999;
    defparam sub_2065_add_2_17.INJECT1_0 = "NO";
    defparam sub_2065_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26673), .COUT(n26674));
    defparam sub_2065_add_2_15.INIT0 = 16'h5999;
    defparam sub_2065_add_2_15.INIT1 = 16'h5999;
    defparam sub_2065_add_2_15.INJECT1_0 = "NO";
    defparam sub_2065_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26672), .COUT(n26673));
    defparam sub_2065_add_2_13.INIT0 = 16'h5999;
    defparam sub_2065_add_2_13.INIT1 = 16'h5999;
    defparam sub_2065_add_2_13.INJECT1_0 = "NO";
    defparam sub_2065_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26671), .COUT(n26672));
    defparam sub_2065_add_2_11.INIT0 = 16'h5999;
    defparam sub_2065_add_2_11.INIT1 = 16'h5999;
    defparam sub_2065_add_2_11.INJECT1_0 = "NO";
    defparam sub_2065_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26670), .COUT(n26671));
    defparam sub_2065_add_2_9.INIT0 = 16'h5999;
    defparam sub_2065_add_2_9.INIT1 = 16'h5999;
    defparam sub_2065_add_2_9.INJECT1_0 = "NO";
    defparam sub_2065_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26669), .COUT(n26670));
    defparam sub_2065_add_2_7.INIT0 = 16'h5999;
    defparam sub_2065_add_2_7.INIT1 = 16'h5999;
    defparam sub_2065_add_2_7.INJECT1_0 = "NO";
    defparam sub_2065_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26668), .COUT(n26669));
    defparam sub_2065_add_2_5.INIT0 = 16'h5999;
    defparam sub_2065_add_2_5.INIT1 = 16'h5999;
    defparam sub_2065_add_2_5.INJECT1_0 = "NO";
    defparam sub_2065_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26667), .COUT(n26668));
    defparam sub_2065_add_2_3.INIT0 = 16'h5999;
    defparam sub_2065_add_2_3.INIT1 = 16'h5999;
    defparam sub_2065_add_2_3.INJECT1_0 = "NO";
    defparam sub_2065_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26667));
    defparam sub_2065_add_2_1.INIT0 = 16'h0000;
    defparam sub_2065_add_2_1.INIT1 = 16'h5999;
    defparam sub_2065_add_2_1.INJECT1_0 = "NO";
    defparam sub_2065_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26666), .S1(n8089));
    defparam sub_2066_add_2_33.INIT0 = 16'hf555;
    defparam sub_2066_add_2_33.INIT1 = 16'h0000;
    defparam sub_2066_add_2_33.INJECT1_0 = "NO";
    defparam sub_2066_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26665), .COUT(n26666));
    defparam sub_2066_add_2_31.INIT0 = 16'hf555;
    defparam sub_2066_add_2_31.INIT1 = 16'hf555;
    defparam sub_2066_add_2_31.INJECT1_0 = "NO";
    defparam sub_2066_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26664), .COUT(n26665));
    defparam sub_2066_add_2_29.INIT0 = 16'hf555;
    defparam sub_2066_add_2_29.INIT1 = 16'hf555;
    defparam sub_2066_add_2_29.INJECT1_0 = "NO";
    defparam sub_2066_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26663), .COUT(n26664));
    defparam sub_2066_add_2_27.INIT0 = 16'hf555;
    defparam sub_2066_add_2_27.INIT1 = 16'hf555;
    defparam sub_2066_add_2_27.INJECT1_0 = "NO";
    defparam sub_2066_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26662), .COUT(n26663));
    defparam sub_2066_add_2_25.INIT0 = 16'hf555;
    defparam sub_2066_add_2_25.INIT1 = 16'hf555;
    defparam sub_2066_add_2_25.INJECT1_0 = "NO";
    defparam sub_2066_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26661), .COUT(n26662));
    defparam sub_2066_add_2_23.INIT0 = 16'hf555;
    defparam sub_2066_add_2_23.INIT1 = 16'hf555;
    defparam sub_2066_add_2_23.INJECT1_0 = "NO";
    defparam sub_2066_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26660), .COUT(n26661));
    defparam sub_2066_add_2_21.INIT0 = 16'hf555;
    defparam sub_2066_add_2_21.INIT1 = 16'hf555;
    defparam sub_2066_add_2_21.INJECT1_0 = "NO";
    defparam sub_2066_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26659), .COUT(n26660));
    defparam sub_2066_add_2_19.INIT0 = 16'hf555;
    defparam sub_2066_add_2_19.INIT1 = 16'hf555;
    defparam sub_2066_add_2_19.INJECT1_0 = "NO";
    defparam sub_2066_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26658), .COUT(n26659));
    defparam sub_2066_add_2_17.INIT0 = 16'hf555;
    defparam sub_2066_add_2_17.INIT1 = 16'hf555;
    defparam sub_2066_add_2_17.INJECT1_0 = "NO";
    defparam sub_2066_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26657), .COUT(n26658));
    defparam sub_2066_add_2_15.INIT0 = 16'hf555;
    defparam sub_2066_add_2_15.INIT1 = 16'hf555;
    defparam sub_2066_add_2_15.INJECT1_0 = "NO";
    defparam sub_2066_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26656), .COUT(n26657));
    defparam sub_2066_add_2_13.INIT0 = 16'hf555;
    defparam sub_2066_add_2_13.INIT1 = 16'hf555;
    defparam sub_2066_add_2_13.INJECT1_0 = "NO";
    defparam sub_2066_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26655), .COUT(n26656));
    defparam sub_2066_add_2_11.INIT0 = 16'hf555;
    defparam sub_2066_add_2_11.INIT1 = 16'hf555;
    defparam sub_2066_add_2_11.INJECT1_0 = "NO";
    defparam sub_2066_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26654), .COUT(n26655));
    defparam sub_2066_add_2_9.INIT0 = 16'hf555;
    defparam sub_2066_add_2_9.INIT1 = 16'hf555;
    defparam sub_2066_add_2_9.INJECT1_0 = "NO";
    defparam sub_2066_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26653), .COUT(n26654));
    defparam sub_2066_add_2_7.INIT0 = 16'hf555;
    defparam sub_2066_add_2_7.INIT1 = 16'hf555;
    defparam sub_2066_add_2_7.INJECT1_0 = "NO";
    defparam sub_2066_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    CCU2D sub_2066_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26652), .COUT(n26653));
    defparam sub_2066_add_2_5.INIT0 = 16'hf555;
    defparam sub_2066_add_2_5.INIT1 = 16'hf555;
    defparam sub_2066_add_2_5.INJECT1_0 = "NO";
    defparam sub_2066_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26651), .COUT(n26652));
    defparam sub_2066_add_2_3.INIT0 = 16'hf555;
    defparam sub_2066_add_2_3.INIT1 = 16'hf555;
    defparam sub_2066_add_2_3.INJECT1_0 = "NO";
    defparam sub_2066_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26651));
    defparam sub_2066_add_2_1.INIT0 = 16'h0000;
    defparam sub_2066_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2066_add_2_1.INJECT1_0 = "NO";
    defparam sub_2066_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31408), .PD(n17034), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1S3IX count_2673__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i1.GSR = "ENABLED";
    FD1S3IX count_2673__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i2.GSR = "ENABLED";
    FD1S3IX count_2673__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i3.GSR = "ENABLED";
    FD1S3IX count_2673__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i4.GSR = "ENABLED";
    FD1S3IX count_2673__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i5.GSR = "ENABLED";
    FD1S3IX count_2673__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i6.GSR = "ENABLED";
    FD1S3IX count_2673__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i7.GSR = "ENABLED";
    FD1S3IX count_2673__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i8.GSR = "ENABLED";
    FD1S3IX count_2673__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i9.GSR = "ENABLED";
    FD1S3IX count_2673__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i10.GSR = "ENABLED";
    FD1S3IX count_2673__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i11.GSR = "ENABLED";
    FD1S3IX count_2673__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i12.GSR = "ENABLED";
    FD1S3IX count_2673__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i13.GSR = "ENABLED";
    FD1S3IX count_2673__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i14.GSR = "ENABLED";
    FD1S3IX count_2673__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i15.GSR = "ENABLED";
    FD1S3IX count_2673__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i16.GSR = "ENABLED";
    FD1S3IX count_2673__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i17.GSR = "ENABLED";
    FD1S3IX count_2673__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i18.GSR = "ENABLED";
    FD1S3IX count_2673__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i19.GSR = "ENABLED";
    FD1S3IX count_2673__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i20.GSR = "ENABLED";
    FD1S3IX count_2673__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i21.GSR = "ENABLED";
    FD1S3IX count_2673__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i22.GSR = "ENABLED";
    FD1S3IX count_2673__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i23.GSR = "ENABLED";
    FD1S3IX count_2673__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i24.GSR = "ENABLED";
    FD1S3IX count_2673__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i25.GSR = "ENABLED";
    FD1S3IX count_2673__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i26.GSR = "ENABLED";
    FD1S3IX count_2673__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i27.GSR = "ENABLED";
    FD1S3IX count_2673__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i28.GSR = "ENABLED";
    FD1S3IX count_2673__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i29.GSR = "ENABLED";
    FD1S3IX count_2673__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i30.GSR = "ENABLED";
    FD1S3IX count_2673__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31408), .CD(n17034), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D count_2673_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27002), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_33.INIT1 = 16'h0000;
    defparam count_2673_add_4_33.INJECT1_0 = "NO";
    defparam count_2673_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27001), .COUT(n27002), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_31.INJECT1_0 = "NO";
    defparam count_2673_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27000), .COUT(n27001), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_29.INJECT1_0 = "NO";
    defparam count_2673_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26999), .COUT(n27000), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_27.INJECT1_0 = "NO";
    defparam count_2673_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26998), .COUT(n26999), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_25.INJECT1_0 = "NO";
    defparam count_2673_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26997), .COUT(n26998), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_23.INJECT1_0 = "NO";
    defparam count_2673_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26996), .COUT(n26997), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2673_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_21.INJECT1_0 = "NO";
    defparam count_2673_add_4_21.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module EncoderPeripheral
//

module EncoderPeripheral (\register_addr[0] , n31431, prev_select, debug_c_c, 
            n31470, \read_size[0] , n15086, n6, encoder_rb_c, encoder_ra_c, 
            read_value, \read_size[2] , n31540, encoder_ri_c, qreset, 
            VCC_net, GND_net, \quadA_delayed[1] , n13938, n6_adj_4, 
            \quadB_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[0] ;
    input n31431;
    output prev_select;
    input debug_c_c;
    input n31470;
    output \read_size[0] ;
    input n15086;
    input n6;
    input encoder_rb_c;
    input encoder_ra_c;
    output [31:0]read_value;
    output \read_size[2] ;
    input n31540;
    input encoder_ri_c;
    input qreset;
    input VCC_net;
    input GND_net;
    output \quadA_delayed[1] ;
    input n13938;
    output n6_adj_4;
    output \quadB_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    wire n29085, n29080, n29105, n29102, n29091, n29084, n29088, 
        n29094, n29104, n29081, n29092, n29093, n29095, n29096, 
        n29082, n29083, n29090, n29098, n29106, n29099, n29086, 
        n29107, n29089, n29108, n29100, n29097, n29087, n29101, 
        n29103;
    wire [31:0]n180;
    
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [4]), 
         .Z(n29085)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_4 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [5]), 
         .Z(n29080)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_4.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_5 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [6]), 
         .Z(n29105)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_5.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_6 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [7]), 
         .Z(n29102)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_6.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_7 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [8]), 
         .Z(n29091)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_7.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_8 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [9]), 
         .Z(n29084)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_8.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_9 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [10]), 
         .Z(n29088)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_9.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_10 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [11]), 
         .Z(n29094)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_10.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_11 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [12]), 
         .Z(n29104)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_11.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_12 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [13]), 
         .Z(n29081)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_12.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_13 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [14]), 
         .Z(n29092)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_13.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_14 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [15]), 
         .Z(n29093)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_14.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_15 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [16]), 
         .Z(n29095)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_15.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_16 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [17]), 
         .Z(n29096)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_16.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_17 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [18]), 
         .Z(n29082)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_17.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_18 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [19]), 
         .Z(n29083)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_18.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_19 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [20]), 
         .Z(n29090)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_19.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_20 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [21]), 
         .Z(n29098)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_20.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_21 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [22]), 
         .Z(n29106)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_21.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_22 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [23]), 
         .Z(n29099)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_22.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_23 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [24]), 
         .Z(n29086)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_23.init = 16'h2020;
    FD1S3AX prev_select_126 (.D(n31470), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam prev_select_126.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_24 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [25]), 
         .Z(n29107)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_24.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_25 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [26]), 
         .Z(n29089)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_25.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_26 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [27]), 
         .Z(n29108)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_26.init = 16'h2020;
    FD1P3IX read_size__i1 (.D(n6), .SP(n15086), .CD(n31431), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_27 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [28]), 
         .Z(n29100)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_27.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_28 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [29]), 
         .Z(n29097)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_28.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_29 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [30]), 
         .Z(n29087)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_29.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_30 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [31]), 
         .Z(n29101)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_30.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_31 (.A(\register_addr[0] ), .B(n31431), .C(\register[1] [0]), 
         .Z(n29103)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_31.init = 16'h2020;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_rb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n180[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_ra_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n180[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i1 (.D(n180[1]), .SP(n15086), .CD(n31431), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_size__i2 (.D(n31540), .SP(n15086), .CD(n31431), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n180[2]), .SP(n15086), .CD(n31431), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n180[3]), .SP(n15086), .CD(n31431), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29085), .SP(n15086), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29080), .SP(n15086), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29105), .SP(n15086), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29102), .SP(n15086), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29091), .SP(n15086), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29084), .SP(n15086), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29088), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29094), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29104), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29081), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29092), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29093), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29095), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29096), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29082), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29083), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29090), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29098), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29106), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29099), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29086), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29107), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29089), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29108), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29100), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29097), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29087), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n29101), .SP(n15086), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i0 (.D(n29103), .SP(n15086), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=680, LSE_RLINE=690 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_ri_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n180[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    QuadratureDecoder q (.\register[1] ({\register[1] }), .debug_c_c(debug_c_c), 
            .qreset(qreset), .VCC_net(VCC_net), .GND_net(GND_net), .encoder_rb_c(encoder_rb_c), 
            .encoder_ra_c(encoder_ra_c), .\quadA_delayed[1] (\quadA_delayed[1] ), 
            .n13938(n13938), .n6(n6_adj_4), .\quadB_delayed[1] (\quadB_delayed[1] )) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(92[20] 96[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder
//

module QuadratureDecoder (\register[1] , debug_c_c, qreset, VCC_net, 
            GND_net, encoder_rb_c, encoder_ra_c, \quadA_delayed[1] , 
            n13938, n6, \quadB_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[1] ;
    input debug_c_c;
    input qreset;
    input VCC_net;
    input GND_net;
    input encoder_rb_c;
    input encoder_ra_c;
    output \quadA_delayed[1] ;
    input n13938;
    output n6;
    output \quadB_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n26521;
    wire [31:0]n4423;
    
    wire n26520, n26519, n26518, n26517, n26516, n26515, n26514, 
        n26513, n26512, n26511, n26510, n26509, n26508, n26507, 
        n26506;
    
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_rb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_ra_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    CCU2D add_1717_33 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n26521), .S0(n4423[30]), 
          .S1(n4423[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_33.INIT0 = 16'h6969;
    defparam add_1717_33.INIT1 = 16'h6969;
    defparam add_1717_33.INJECT1_0 = "NO";
    defparam add_1717_33.INJECT1_1 = "NO";
    CCU2D add_1717_31 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n26520), .COUT(n26521), 
          .S0(n4423[28]), .S1(n4423[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_31.INIT0 = 16'h6969;
    defparam add_1717_31.INIT1 = 16'h6969;
    defparam add_1717_31.INJECT1_0 = "NO";
    defparam add_1717_31.INJECT1_1 = "NO";
    CCU2D add_1717_29 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n26519), .COUT(n26520), 
          .S0(n4423[26]), .S1(n4423[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_29.INIT0 = 16'h6969;
    defparam add_1717_29.INIT1 = 16'h6969;
    defparam add_1717_29.INJECT1_0 = "NO";
    defparam add_1717_29.INJECT1_1 = "NO";
    CCU2D add_1717_27 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n26518), .COUT(n26519), 
          .S0(n4423[24]), .S1(n4423[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_27.INIT0 = 16'h6969;
    defparam add_1717_27.INIT1 = 16'h6969;
    defparam add_1717_27.INJECT1_0 = "NO";
    defparam add_1717_27.INJECT1_1 = "NO";
    CCU2D add_1717_25 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n26517), .COUT(n26518), 
          .S0(n4423[22]), .S1(n4423[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_25.INIT0 = 16'h6969;
    defparam add_1717_25.INIT1 = 16'h6969;
    defparam add_1717_25.INJECT1_0 = "NO";
    defparam add_1717_25.INJECT1_1 = "NO";
    CCU2D add_1717_23 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n26516), .COUT(n26517), 
          .S0(n4423[20]), .S1(n4423[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_23.INIT0 = 16'h6969;
    defparam add_1717_23.INIT1 = 16'h6969;
    defparam add_1717_23.INJECT1_0 = "NO";
    defparam add_1717_23.INJECT1_1 = "NO";
    CCU2D add_1717_21 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n26515), .COUT(n26516), 
          .S0(n4423[18]), .S1(n4423[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_21.INIT0 = 16'h6969;
    defparam add_1717_21.INIT1 = 16'h6969;
    defparam add_1717_21.INJECT1_0 = "NO";
    defparam add_1717_21.INJECT1_1 = "NO";
    CCU2D add_1717_19 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n26514), .COUT(n26515), 
          .S0(n4423[16]), .S1(n4423[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_19.INIT0 = 16'h6969;
    defparam add_1717_19.INIT1 = 16'h6969;
    defparam add_1717_19.INJECT1_0 = "NO";
    defparam add_1717_19.INJECT1_1 = "NO";
    CCU2D add_1717_17 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n26513), .COUT(n26514), 
          .S0(n4423[14]), .S1(n4423[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_17.INIT0 = 16'h6969;
    defparam add_1717_17.INIT1 = 16'h6969;
    defparam add_1717_17.INJECT1_0 = "NO";
    defparam add_1717_17.INJECT1_1 = "NO";
    CCU2D add_1717_15 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n26512), .COUT(n26513), 
          .S0(n4423[12]), .S1(n4423[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_15.INIT0 = 16'h6969;
    defparam add_1717_15.INIT1 = 16'h6969;
    defparam add_1717_15.INJECT1_0 = "NO";
    defparam add_1717_15.INJECT1_1 = "NO";
    CCU2D add_1717_13 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n26511), .COUT(n26512), 
          .S0(n4423[10]), .S1(n4423[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_13.INIT0 = 16'h6969;
    defparam add_1717_13.INIT1 = 16'h6969;
    defparam add_1717_13.INJECT1_0 = "NO";
    defparam add_1717_13.INJECT1_1 = "NO";
    CCU2D add_1717_11 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n26510), .COUT(n26511), 
          .S0(n4423[8]), .S1(n4423[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_11.INIT0 = 16'h6969;
    defparam add_1717_11.INIT1 = 16'h6969;
    defparam add_1717_11.INJECT1_0 = "NO";
    defparam add_1717_11.INJECT1_1 = "NO";
    CCU2D add_1717_9 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n26509), .COUT(n26510), 
          .S0(n4423[6]), .S1(n4423[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_9.INIT0 = 16'h6969;
    defparam add_1717_9.INIT1 = 16'h6969;
    defparam add_1717_9.INJECT1_0 = "NO";
    defparam add_1717_9.INJECT1_1 = "NO";
    CCU2D add_1717_7 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n26508), .COUT(n26509), 
          .S0(n4423[4]), .S1(n4423[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_7.INIT0 = 16'h6969;
    defparam add_1717_7.INIT1 = 16'h6969;
    defparam add_1717_7.INJECT1_0 = "NO";
    defparam add_1717_7.INJECT1_1 = "NO";
    CCU2D add_1717_5 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n26507), .COUT(n26508), 
          .S0(n4423[2]), .S1(n4423[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_5.INIT0 = 16'h6969;
    defparam add_1717_5.INIT1 = 16'h6969;
    defparam add_1717_5.INJECT1_0 = "NO";
    defparam add_1717_5.INJECT1_1 = "NO";
    CCU2D add_1717_3 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n26506), .COUT(n26507), 
          .S0(n4423[0]), .S1(n4423[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_3.INIT0 = 16'h9696;
    defparam add_1717_3.INIT1 = 16'h6969;
    defparam add_1717_3.INJECT1_0 = "NO";
    defparam add_1717_3.INJECT1_1 = "NO";
    CCU2D add_1717_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26506));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1717_1.INIT0 = 16'hF000;
    defparam add_1717_1.INIT1 = 16'h6666;
    defparam add_1717_1.INJECT1_0 = "NO";
    defparam add_1717_1.INJECT1_1 = "NO";
    FD1P3IX count__i31 (.D(n4423[31]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4423[30]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n4423[29]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n4423[28]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n4423[27]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n4423[26]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n4423[25]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n4423[24]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n4423[23]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n4423[22]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n4423[21]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n4423[20]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n4423[19]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n4423[18]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n4423[17]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n4423[16]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n4423[15]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n4423[14]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n4423[13]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n4423[12]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n4423[11]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n4423[10]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n4423[9]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n4423[8]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n4423[7]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n4423[6]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n4423[5]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n4423[4]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n4423[3]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n4423[2]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n4423[1]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    FD1P3IX count__i0 (.D(n4423[0]), .SP(n13938), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed[0]), .CK(debug_c_c), .Q(\quadA_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(\quadA_delayed[1] ), .CK(debug_c_c), .Q(quadA_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP_SP(factor=120000) 
//

module \ClockDividerP_SP(factor=120000)  (n29791, debug_c_0, debug_c_c, 
            n31511, n2860, GND_net) /* synthesis syn_module_defined=1 */ ;
    output n29791;
    output debug_c_0;
    input debug_c_c;
    input n31511;
    input n2860;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(86[13:18])
    
    wire n21, n19, n25, n38, n34, n26, n31480, n20, n36, n30, 
        n32, n22, n29535, n29679, n29533, n29661, n29541, n27788;
    wire [31:0]n134;
    
    wire n26938, n26937, n26936, n26935, n26934, n26933, n26932, 
        n26931, n26930, n26929, n26928, n26927, n26926, n26925, 
        n26924, n26923;
    
    LUT4 i9_4_lut (.A(count[5]), .B(count[16]), .C(count[12]), .D(count[14]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(count[7]), .B(count[15]), .C(count[4]), .D(count[10]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut_rep_337 (.A(n25), .B(n38), .C(n34), .D(n26), .Z(n31480)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i19_4_lut_rep_337.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[1]), .B(count[0]), .C(count[2]), .D(count[3]), 
         .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[11]), .B(count[13]), .Z(n25)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(count[6]), .B(n36), .C(n30), .D(count[9]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(count[20]), .B(count[31]), .C(count[24]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(count[21]), .B(count[17]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i16_4_lut (.A(count[26]), .B(n32), .C(n22), .D(count[29]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(count[18]), .B(count[28]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(count[25]), .B(count[23]), .C(count[8]), .D(count[27]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[19]), .B(count[22]), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i22331_4_lut (.A(n31480), .B(n29535), .C(n29679), .D(n29533), 
         .Z(n29791)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i22331_4_lut.init = 16'h4000;
    LUT4 i21981_2_lut (.A(count[10]), .B(count[12]), .Z(n29535)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21981_2_lut.init = 16'h8888;
    LUT4 i22119_4_lut (.A(count[3]), .B(n29661), .C(n29541), .D(count[0]), 
         .Z(n29679)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22119_4_lut.init = 16'h8000;
    LUT4 i21979_2_lut (.A(count[2]), .B(count[5]), .Z(n29533)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21979_2_lut.init = 16'h8888;
    LUT4 i22101_4_lut (.A(count[1]), .B(count[16]), .C(count[4]), .D(count[15]), 
         .Z(n29661)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22101_4_lut.init = 16'h8000;
    LUT4 i21987_2_lut (.A(count[7]), .B(count[14]), .Z(n29541)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21987_2_lut.init = 16'h8888;
    FD1S3IX clk_o_13 (.D(n27788), .CK(debug_c_c), .CD(n31511), .Q(debug_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(88[9] 107[6])
    defparam clk_o_13.GSR = "ENABLED";
    FD1S3IX count_2671__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2860), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i0.GSR = "ENABLED";
    CCU2D count_2671_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26938), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_33.INIT1 = 16'h0000;
    defparam count_2671_add_4_33.INJECT1_0 = "NO";
    defparam count_2671_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26937), .COUT(n26938), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_31.INJECT1_0 = "NO";
    defparam count_2671_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26936), .COUT(n26937), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_29.INJECT1_0 = "NO";
    defparam count_2671_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26935), .COUT(n26936), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_27.INJECT1_0 = "NO";
    defparam count_2671_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26934), .COUT(n26935), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_25.INJECT1_0 = "NO";
    defparam count_2671_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26933), .COUT(n26934), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_23.INJECT1_0 = "NO";
    defparam count_2671_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26932), .COUT(n26933), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_21.INJECT1_0 = "NO";
    defparam count_2671_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26931), .COUT(n26932), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_19.INJECT1_0 = "NO";
    defparam count_2671_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26930), .COUT(n26931), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_17.INJECT1_0 = "NO";
    defparam count_2671_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26929), .COUT(n26930), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_15.INJECT1_0 = "NO";
    defparam count_2671_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26928), .COUT(n26929), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_13.INJECT1_0 = "NO";
    defparam count_2671_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26927), .COUT(n26928), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_11.INJECT1_0 = "NO";
    defparam count_2671_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26926), .COUT(n26927), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_9.INJECT1_0 = "NO";
    defparam count_2671_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26925), .COUT(n26926), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_7.INJECT1_0 = "NO";
    defparam count_2671_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26924), .COUT(n26925), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_5.INJECT1_0 = "NO";
    defparam count_2671_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26923), .COUT(n26924), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_3.INJECT1_0 = "NO";
    defparam count_2671_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26923), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671_add_4_1.INIT0 = 16'hF000;
    defparam count_2671_add_4_1.INIT1 = 16'h0555;
    defparam count_2671_add_4_1.INJECT1_0 = "NO";
    defparam count_2671_add_4_1.INJECT1_1 = "NO";
    LUT4 i22375_4_lut_4_lut (.A(n31480), .B(n20), .C(n19), .D(n21), 
         .Z(n27788)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i22375_4_lut_4_lut.init = 16'h0001;
    FD1S3IX count_2671__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2860), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i1.GSR = "ENABLED";
    FD1S3IX count_2671__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2860), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i2.GSR = "ENABLED";
    FD1S3IX count_2671__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2860), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i3.GSR = "ENABLED";
    FD1S3IX count_2671__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2860), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i4.GSR = "ENABLED";
    FD1S3IX count_2671__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2860), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i5.GSR = "ENABLED";
    FD1S3IX count_2671__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2860), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i6.GSR = "ENABLED";
    FD1S3IX count_2671__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2860), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i7.GSR = "ENABLED";
    FD1S3IX count_2671__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2860), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i8.GSR = "ENABLED";
    FD1S3IX count_2671__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2860), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i9.GSR = "ENABLED";
    FD1S3IX count_2671__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i10.GSR = "ENABLED";
    FD1S3IX count_2671__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i11.GSR = "ENABLED";
    FD1S3IX count_2671__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i12.GSR = "ENABLED";
    FD1S3IX count_2671__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i13.GSR = "ENABLED";
    FD1S3IX count_2671__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i14.GSR = "ENABLED";
    FD1S3IX count_2671__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i15.GSR = "ENABLED";
    FD1S3IX count_2671__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i16.GSR = "ENABLED";
    FD1S3IX count_2671__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i17.GSR = "ENABLED";
    FD1S3IX count_2671__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i18.GSR = "ENABLED";
    FD1S3IX count_2671__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i19.GSR = "ENABLED";
    FD1S3IX count_2671__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i20.GSR = "ENABLED";
    FD1S3IX count_2671__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i21.GSR = "ENABLED";
    FD1S3IX count_2671__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i22.GSR = "ENABLED";
    FD1S3IX count_2671__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i23.GSR = "ENABLED";
    FD1S3IX count_2671__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i24.GSR = "ENABLED";
    FD1S3IX count_2671__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i25.GSR = "ENABLED";
    FD1S3IX count_2671__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i26.GSR = "ENABLED";
    FD1S3IX count_2671__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i27.GSR = "ENABLED";
    FD1S3IX count_2671__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i28.GSR = "ENABLED";
    FD1S3IX count_2671__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i29.GSR = "ENABLED";
    FD1S3IX count_2671__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i30.GSR = "ENABLED";
    FD1S3IX count_2671__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2860), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2671__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module EncoderPeripheral_U11
//

module EncoderPeripheral_U11 (\read_size[0] , debug_c_c, n14145, n31426, 
            n31449, prev_select, n31464, \read_size[2] , n31477, read_value, 
            \register_addr[0] , encoder_la_c, encoder_lb_c, n59, n57, 
            n45, \quadA_delayed[1] , qreset, n6, \quadB_delayed[1] , 
            n13938, n97, encoder_li_c, GND_net, \register[1][0] , 
            VCC_net, \register[1][19] , \register[1][20] , \register[1][26] ) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n14145;
    input n31426;
    input n31449;
    output prev_select;
    input n31464;
    output \read_size[2] ;
    input n31477;
    output [31:0]read_value;
    input \register_addr[0] ;
    input encoder_la_c;
    input encoder_lb_c;
    input n59;
    input n57;
    input n45;
    input \quadA_delayed[1] ;
    input qreset;
    input n6;
    input \quadB_delayed[1] ;
    output n13938;
    input n97;
    input encoder_li_c;
    input GND_net;
    output \register[1][0] ;
    input VCC_net;
    output \register[1][19] ;
    output \register[1][20] ;
    output \register[1][26] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]n100;
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n6_adj_19;
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n15144;
    
    FD1P3IX read_size__i1 (.D(n31449), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3AX prev_select_126 (.D(n31464), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam prev_select_126.GSR = "ENABLED";
    FD1P3IX read_size__i2 (.D(n31477), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i28.GSR = "ENABLED";
    LUT4 i15001_2_lut (.A(\register[1] [31]), .B(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15001_2_lut.init = 16'h8888;
    LUT4 i15002_2_lut (.A(\register[1] [30]), .B(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15002_2_lut.init = 16'h8888;
    LUT4 i15003_2_lut (.A(\register[1] [29]), .B(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15003_2_lut.init = 16'h8888;
    LUT4 i15006_2_lut (.A(\register[1] [28]), .B(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15006_2_lut.init = 16'h8888;
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n100[2]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n100[1]), .SP(n14145), .CD(n31426), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i15007_2_lut (.A(\register[1] [27]), .B(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15007_2_lut.init = 16'h8888;
    LUT4 i15008_2_lut (.A(\register[1] [25]), .B(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15008_2_lut.init = 16'h8888;
    LUT4 i15009_2_lut (.A(\register[1] [24]), .B(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15009_2_lut.init = 16'h8888;
    LUT4 i15010_2_lut (.A(\register[1] [23]), .B(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15010_2_lut.init = 16'h8888;
    LUT4 i15011_2_lut (.A(\register[1] [22]), .B(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15011_2_lut.init = 16'h8888;
    LUT4 i15012_2_lut (.A(\register[1] [21]), .B(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15012_2_lut.init = 16'h8888;
    LUT4 i15013_2_lut (.A(\register[1] [18]), .B(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15013_2_lut.init = 16'h8888;
    LUT4 i15014_2_lut (.A(\register[1] [17]), .B(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15014_2_lut.init = 16'h8888;
    LUT4 i15015_2_lut (.A(\register[1] [16]), .B(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15015_2_lut.init = 16'h8888;
    LUT4 i15016_2_lut (.A(\register[1] [15]), .B(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15016_2_lut.init = 16'h8888;
    LUT4 i15017_2_lut (.A(\register[1] [14]), .B(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15017_2_lut.init = 16'h8888;
    LUT4 i15018_2_lut (.A(\register[1] [13]), .B(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15018_2_lut.init = 16'h8888;
    LUT4 i15019_2_lut (.A(\register[1] [12]), .B(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15019_2_lut.init = 16'h8888;
    LUT4 i15020_2_lut (.A(\register[1] [11]), .B(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15020_2_lut.init = 16'h8888;
    LUT4 i15021_2_lut (.A(\register[1] [10]), .B(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15021_2_lut.init = 16'h8888;
    LUT4 i15022_2_lut (.A(\register[1] [9]), .B(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15022_2_lut.init = 16'h8888;
    LUT4 i15023_2_lut (.A(\register[1] [8]), .B(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15023_2_lut.init = 16'h8888;
    LUT4 i15024_2_lut (.A(\register[1] [7]), .B(\register_addr[0] ), .Z(n100[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15024_2_lut.init = 16'h8888;
    LUT4 i15025_2_lut (.A(\register[1] [6]), .B(\register_addr[0] ), .Z(n100[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15025_2_lut.init = 16'h8888;
    LUT4 i15026_2_lut (.A(\register[1] [5]), .B(\register_addr[0] ), .Z(n100[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15026_2_lut.init = 16'h8888;
    LUT4 i15027_2_lut (.A(\register[1] [4]), .B(\register_addr[0] ), .Z(n100[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15027_2_lut.init = 16'h8888;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_la_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n100[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_lb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n100[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i19 (.D(n59), .SP(n14145), .CK(debug_c_c), .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n57), .SP(n14145), .CK(debug_c_c), .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n45), .SP(n14145), .CK(debug_c_c), .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i26.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(\quadA_delayed[1] ), .B(qreset), .C(n6), .D(\quadB_delayed[1] ), 
         .Z(n13938)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(62[18:35])
    defparam i1_4_lut.init = 16'hedde;
    FD1P3AX read_value__i0 (.D(n97), .SP(n14145), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=669, LSE_RLINE=679 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_li_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n100[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_3 (.A(quadA_delayed[1]), .B(qreset), .C(n6_adj_19), 
         .D(quadB_delayed[1]), .Z(n15144)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(62[18:35])
    defparam i1_4_lut_adj_3.init = 16'hedde;
    QuadratureDecoder_U6 q (.GND_net(GND_net), .quadA_delayed({Open_2, quadA_delayed[1], 
            Open_3}), .\register[1] ({\register[1] [31:27], \register[1][26] , 
            \register[1] [25:21], \register[1][20] , \register[1][19] , 
            \register[1] [18:1], \register[1][0] }), .debug_c_c(debug_c_c), 
            .qreset(qreset), .VCC_net(VCC_net), .encoder_lb_c(encoder_lb_c), 
            .n15144(n15144), .encoder_la_c(encoder_la_c), .\quadB_delayed[1] (quadB_delayed[1]), 
            .n6(n6_adj_19)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(92[20] 96[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder_U6
//

module QuadratureDecoder_U6 (GND_net, quadA_delayed, \register[1] , debug_c_c, 
            qreset, VCC_net, encoder_lb_c, n15144, encoder_la_c, \quadB_delayed[1] , 
            n6) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [2:0]quadA_delayed;
    output [31:0]\register[1] ;
    input debug_c_c;
    input qreset;
    input VCC_net;
    input encoder_lb_c;
    input n15144;
    input encoder_la_c;
    output \quadB_delayed[1] ;
    output n6;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n26438;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [31:0]n4357;
    wire [2:0]quadA_delayed_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n26453, n26452;
    wire [31:0]n100;
    
    wire n26451, n26450, n26449, n26448, n26447, n26446, n26445, 
        n26444, n26443, n26442, n26441, n26440, n26439;
    
    CCU2D add_1683_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26438));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_1.INIT0 = 16'hF000;
    defparam add_1683_1.INIT1 = 16'h6666;
    defparam add_1683_1.INJECT1_0 = "NO";
    defparam add_1683_1.INJECT1_1 = "NO";
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_lb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    FD1P3IX count__i0 (.D(n4357[0]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_la_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed_c[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    CCU2D add_1683_33 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n26453), .S0(n4357[30]), 
          .S1(n4357[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_33.INIT0 = 16'h6969;
    defparam add_1683_33.INIT1 = 16'h6969;
    defparam add_1683_33.INJECT1_0 = "NO";
    defparam add_1683_33.INJECT1_1 = "NO";
    CCU2D add_1683_31 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n26452), .COUT(n26453), 
          .S0(n100[28]), .S1(n100[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_31.INIT0 = 16'h6969;
    defparam add_1683_31.INIT1 = 16'h6969;
    defparam add_1683_31.INJECT1_0 = "NO";
    defparam add_1683_31.INJECT1_1 = "NO";
    CCU2D add_1683_29 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n26451), .COUT(n26452), 
          .S0(n100[26]), .S1(n100[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_29.INIT0 = 16'h6969;
    defparam add_1683_29.INIT1 = 16'h6969;
    defparam add_1683_29.INJECT1_0 = "NO";
    defparam add_1683_29.INJECT1_1 = "NO";
    CCU2D add_1683_27 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n26450), .COUT(n26451), 
          .S0(n100[24]), .S1(n100[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_27.INIT0 = 16'h6969;
    defparam add_1683_27.INIT1 = 16'h6969;
    defparam add_1683_27.INJECT1_0 = "NO";
    defparam add_1683_27.INJECT1_1 = "NO";
    CCU2D add_1683_25 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n26449), .COUT(n26450), 
          .S0(n100[22]), .S1(n100[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_25.INIT0 = 16'h6969;
    defparam add_1683_25.INIT1 = 16'h6969;
    defparam add_1683_25.INJECT1_0 = "NO";
    defparam add_1683_25.INJECT1_1 = "NO";
    FD1P3IX count__i31 (.D(n4357[31]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4357[30]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    CCU2D add_1683_23 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n26448), .COUT(n26449), 
          .S0(n100[20]), .S1(n100[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_23.INIT0 = 16'h6969;
    defparam add_1683_23.INIT1 = 16'h6969;
    defparam add_1683_23.INJECT1_0 = "NO";
    defparam add_1683_23.INJECT1_1 = "NO";
    CCU2D add_1683_21 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n26447), .COUT(n26448), 
          .S0(n100[18]), .S1(n100[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_21.INIT0 = 16'h6969;
    defparam add_1683_21.INIT1 = 16'h6969;
    defparam add_1683_21.INJECT1_0 = "NO";
    defparam add_1683_21.INJECT1_1 = "NO";
    CCU2D add_1683_19 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n26446), .COUT(n26447), 
          .S0(n100[16]), .S1(n100[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_19.INIT0 = 16'h6969;
    defparam add_1683_19.INIT1 = 16'h6969;
    defparam add_1683_19.INJECT1_0 = "NO";
    defparam add_1683_19.INJECT1_1 = "NO";
    CCU2D add_1683_17 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n26445), .COUT(n26446), 
          .S0(n100[14]), .S1(n100[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_17.INIT0 = 16'h6969;
    defparam add_1683_17.INIT1 = 16'h6969;
    defparam add_1683_17.INJECT1_0 = "NO";
    defparam add_1683_17.INJECT1_1 = "NO";
    CCU2D add_1683_15 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n26444), .COUT(n26445), 
          .S0(n100[12]), .S1(n100[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_15.INIT0 = 16'h6969;
    defparam add_1683_15.INIT1 = 16'h6969;
    defparam add_1683_15.INJECT1_0 = "NO";
    defparam add_1683_15.INJECT1_1 = "NO";
    CCU2D add_1683_13 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n26443), .COUT(n26444), 
          .S0(n100[10]), .S1(n100[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_13.INIT0 = 16'h6969;
    defparam add_1683_13.INIT1 = 16'h6969;
    defparam add_1683_13.INJECT1_0 = "NO";
    defparam add_1683_13.INJECT1_1 = "NO";
    CCU2D add_1683_11 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n26442), .COUT(n26443), 
          .S0(n100[8]), .S1(n100[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_11.INIT0 = 16'h6969;
    defparam add_1683_11.INIT1 = 16'h6969;
    defparam add_1683_11.INJECT1_0 = "NO";
    defparam add_1683_11.INJECT1_1 = "NO";
    CCU2D add_1683_9 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n26441), .COUT(n26442), 
          .S0(n100[6]), .S1(n100[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_9.INIT0 = 16'h6969;
    defparam add_1683_9.INIT1 = 16'h6969;
    defparam add_1683_9.INJECT1_0 = "NO";
    defparam add_1683_9.INJECT1_1 = "NO";
    CCU2D add_1683_7 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n26440), .COUT(n26441), 
          .S0(n100[4]), .S1(n100[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_7.INIT0 = 16'h6969;
    defparam add_1683_7.INIT1 = 16'h6969;
    defparam add_1683_7.INJECT1_0 = "NO";
    defparam add_1683_7.INJECT1_1 = "NO";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n100[1]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n100[2]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n100[3]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n100[4]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n100[5]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n100[6]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n100[7]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n100[8]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n100[9]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n100[10]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n100[11]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n100[12]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n100[13]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n100[14]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n100[15]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n100[16]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n100[17]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n100[18]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n100[19]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n100[20]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n100[21]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n100[22]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n100[23]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n100[24]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n100[25]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n100[26]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n100[27]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n100[28]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n100[29]), .SP(n15144), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed_c[0]), .CK(debug_c_c), .Q(quadA_delayed[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(quadA_delayed[1]), .CK(debug_c_c), .Q(quadA_delayed_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    CCU2D add_1683_5 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n26439), .COUT(n26440), 
          .S0(n100[2]), .S1(n100[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_5.INIT0 = 16'h6969;
    defparam add_1683_5.INIT1 = 16'h6969;
    defparam add_1683_5.INJECT1_0 = "NO";
    defparam add_1683_5.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed_c[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    CCU2D add_1683_3 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n26438), .COUT(n26439), 
          .S0(n4357[0]), .S1(n100[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_3.INIT0 = 16'h9696;
    defparam add_1683_3.INIT1 = 16'h6969;
    defparam add_1683_3.INJECT1_0 = "NO";
    defparam add_1683_3.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (read_value, debug_c_c, n2857, 
            n31511, n3921, VCC_net, GND_net, Stepper_A_nFault_c, \read_size[0] , 
            n29257, Stepper_A_M0_c_0, databus, limit_latched, prev_limit_latched, 
            n9330, prev_select, n31444, Stepper_A_M1_c_1, \register_addr[0] , 
            \register_addr[1] , n224, n32, n32_adj_1, prev_step_clk, 
            step_clk, n31418, n22, prev_step_clk_adj_2, n34, step_clk_adj_3, 
            n31420, n24, n31427, \register_addr[5] , n31496, n29270, 
            n31575, n27441, \read_size[2] , n29256, Stepper_A_M2_c_2, 
            Stepper_A_Dir_c, Stepper_A_En_c, \control_reg[7] , n12210, 
            Stepper_A_Step_c, limit_c_3, n8653, n31409, n8401, n8367, 
            n16842) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2857;
    input n31511;
    input [31:0]n3921;
    input VCC_net;
    input GND_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n29257;
    output Stepper_A_M0_c_0;
    input [31:0]databus;
    output limit_latched;
    output prev_limit_latched;
    input n9330;
    output prev_select;
    input n31444;
    output Stepper_A_M1_c_1;
    input \register_addr[0] ;
    input \register_addr[1] ;
    output [31:0]n224;
    input n32;
    input n32_adj_1;
    input prev_step_clk;
    input step_clk;
    output n31418;
    output n22;
    input prev_step_clk_adj_2;
    input n34;
    input step_clk_adj_3;
    output n31420;
    output n24;
    input n31427;
    input \register_addr[5] ;
    input n31496;
    input n29270;
    input n31575;
    output n27441;
    output \read_size[2] ;
    input n29256;
    output Stepper_A_M2_c_2;
    output Stepper_A_Dir_c;
    output Stepper_A_En_c;
    output \control_reg[7] ;
    input n12210;
    output Stepper_A_Step_c;
    input limit_c_3;
    input n8653;
    input n31409;
    output n8401;
    output n8367;
    input n16842;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n49, n41, n60, n54, n42, n62, n52, n38, n58, n50, 
        n56, n46, n9555, n29691, fault_latched, n13942, prev_step_clk_c, 
        step_clk_c, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n29698, n29699;
    wire [31:0]n100;
    
    wire n29730, n29700, n26834, n26833, n31416, n22_c, n26832, 
        n26831, n26830, n26829, n26828, n26827, n26826, n26825, 
        n26824, n26823, n26822, n26821, n26820, n26819, n29728, 
        n29729, n29689, n29690;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire int_step;
    wire [7:0]n8652;
    wire [31:0]n7370;
    
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(steps_reg[9]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    FD1P3IX read_value__i0 (.D(n29691), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(steps_reg[3]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[6]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    FD1S3IX steps_reg__i0 (.D(n3921[0]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n29257), .SP(n2857), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n13942), .CD(n31511), 
            .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk_c), .CK(debug_c_c), .Q(prev_step_clk_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31444), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3921[31]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3921[30]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3921[29]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3921[28]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3921[27]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3921[26]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3921[25]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3921[24]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3921[23]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3921[22]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3921[21]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3921[20]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3921[19]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3921[18]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3921[17]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3921[16]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3921[15]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3921[14]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3921[13]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3921[12]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3921[11]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3921[10]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3921[9]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3921[8]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3921[7]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3921[6]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3921[5]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3921[4]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3921[3]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3921[2]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3921[1]), .CK(debug_c_c), .CD(n31511), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i22138_3_lut (.A(Stepper_A_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22138_3_lut.init = 16'hcaca;
    LUT4 i22139_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22139_3_lut.init = 16'hcaca;
    LUT4 i14871_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14871_4_lut.init = 16'hc088;
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i14872_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14872_4_lut.init = 16'hc088;
    LUT4 i14873_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14873_4_lut.init = 16'hc088;
    LUT4 i14874_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14874_4_lut.init = 16'hc088;
    LUT4 i14875_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14875_4_lut.init = 16'hc088;
    LUT4 i14876_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14876_4_lut.init = 16'hc088;
    LUT4 i14877_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14877_4_lut.init = 16'hc088;
    LUT4 i14878_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14878_4_lut.init = 16'hc088;
    LUT4 i14879_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14879_4_lut.init = 16'hc088;
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29730), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29700), .SP(n2857), .CD(n9555), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i14880_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14880_4_lut.init = 16'hc088;
    LUT4 i14881_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14881_4_lut.init = 16'hc088;
    LUT4 i14882_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14882_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26834), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26833), .COUT(n26834), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_273 (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .Z(n31416)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_273.init = 16'h2020;
    LUT4 i14883_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14883_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_4_lut (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .D(n31511), .Z(n22_c)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut.init = 16'h002c;
    LUT4 i14884_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14884_4_lut.init = 16'hc088;
    LUT4 i14885_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14885_4_lut.init = 16'hc088;
    LUT4 i2_3_lut_rep_275 (.A(n32_adj_1), .B(prev_step_clk), .C(step_clk), 
         .Z(n31418)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_275.init = 16'h2020;
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26832), .COUT(n26833), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_adj_1 (.A(n32_adj_1), .B(prev_step_clk), .C(step_clk), 
         .D(n31511), .Z(n22)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_1.init = 16'h002c;
    LUT4 i14886_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14886_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26831), .COUT(n26832), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    LUT4 i14887_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14887_4_lut.init = 16'hc088;
    LUT4 i14888_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14888_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26830), .COUT(n26831), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    LUT4 i14889_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14889_4_lut.init = 16'hc088;
    LUT4 i14890_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14890_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26829), .COUT(n26830), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26828), .COUT(n26829), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    LUT4 i14891_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14891_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26827), .COUT(n26828), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26826), .COUT(n26827), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26825), .COUT(n26826), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26824), .COUT(n26825), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_277 (.A(prev_step_clk_adj_2), .B(n34), .C(step_clk_adj_3), 
         .Z(n31420)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_277.init = 16'h4040;
    LUT4 i14892_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14892_4_lut.init = 16'hc088;
    LUT4 i14893_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14893_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26823), .COUT(n26824), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26822), .COUT(n26823), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 i14894_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14894_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26821), .COUT(n26822), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_adj_2 (.A(prev_step_clk_adj_2), .B(n34), .C(step_clk_adj_3), 
         .D(n31511), .Z(n24)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_2.init = 16'h004a;
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26820), .COUT(n26821), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26819), .COUT(n26820), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk_c), .D1(prev_step_clk_c), 
          .COUT(n26819), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n31427), .B(n31511), .C(\register_addr[5] ), .D(n31496), 
         .Z(n9555)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_4_lut.init = 16'h0222;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31444), .B(prev_select), .C(n29270), 
         .D(n31575), .Z(n13942)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27441)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    PFUMX i22170 (.BLUT(n29728), .ALUT(n29729), .C0(\register_addr[0] ), 
          .Z(n29730));
    FD1P3AX read_size__i2 (.D(n29256), .SP(n2857), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    PFUMX i22131 (.BLUT(n29689), .ALUT(n29690), .C0(\register_addr[1] ), 
          .Z(n29691));
    PFUMX i22140 (.BLUT(n29698), .ALUT(n29699), .C0(\register_addr[1] ), 
          .Z(n29700));
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13942), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13942), .CD(n31511), 
            .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13942), .PD(n31511), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13942), .CD(n31511), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13942), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13942), .PD(n31511), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13942), .CD(n12210), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9330), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9330), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9330), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9330), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9330), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9330), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9330), .PD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9330), .CD(n31511), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=623, LSE_RLINE=636 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i22168_3_lut (.A(Stepper_A_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n29728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22168_3_lut.init = 16'hcaca;
    LUT4 i22169_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n29729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22169_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n31416), .SP(n22_c), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i22129_3_lut (.A(Stepper_A_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n29689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22129_3_lut.init = 16'hcaca;
    LUT4 i14870_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8652[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14870_2_lut.init = 16'h2222;
    LUT4 mux_2001_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7370[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2001_i4_3_lut.init = 16'hcaca;
    LUT4 i14869_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8652[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14869_2_lut.init = 16'h2222;
    LUT4 mux_2001_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7370[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2001_i5_3_lut.init = 16'hcaca;
    LUT4 i14868_2_lut (.A(Stepper_A_Dir_c), .B(\register_addr[0] ), .Z(n8652[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14868_2_lut.init = 16'h2222;
    LUT4 mux_2001_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7370[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2001_i6_3_lut.init = 16'hcaca;
    LUT4 i14867_2_lut (.A(Stepper_A_En_c), .B(\register_addr[0] ), .Z(n8652[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14867_2_lut.init = 16'h2222;
    LUT4 i22130_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n29690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22130_3_lut.init = 16'hcaca;
    LUT4 mux_2001_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7370[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2001_i7_3_lut.init = 16'hcaca;
    LUT4 mux_2001_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n7370[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2001_i8_3_lut.init = 16'hcaca;
    PFUMX mux_2005_i4 (.BLUT(n8652[3]), .ALUT(n7370[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_2005_i5 (.BLUT(n8652[4]), .ALUT(n7370[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_2005_i6 (.BLUT(n8652[5]), .ALUT(n7370[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_2005_i7 (.BLUT(n8652[6]), .ALUT(n7370[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    PFUMX mux_2005_i8 (.BLUT(n8653), .ALUT(n7370[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    ClockDivider_U9 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk_c), 
            .debug_c_c(debug_c_c), .n31511(n31511), .n31409(n31409), .div_factor_reg({div_factor_reg}), 
            .n8401(n8401), .n8367(n8367), .n16842(n16842)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (GND_net, step_clk, debug_c_c, n31511, n31409, 
            div_factor_reg, n8401, n8367, n16842) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31511;
    input n31409;
    input [31:0]div_factor_reg;
    output n8401;
    output n8367;
    input n16842;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26550;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26551, n26549, n26548, n26547, n8332, n26546, n26545, 
        n26544, n26543, n26954;
    wire [31:0]n134;
    
    wire n26953, n26952, n26951, n26950, n26542, n26541, n26949, 
        n26948, n26947, n26946, n26945, n26944, n26943, n26942, 
        n26941, n26940, n26939, n27114, n27113, n27112, n27111, 
        n27110, n27109, n27108, n27107, n27106, n27105, n26540, 
        n27104, n26539, n26538;
    wire [31:0]n40;
    
    wire n26537, n26536, n26535, n26534, n27103, n26533, n26532, 
        n27102, n26531, n26530, n26529, n26528, n26527, n26526, 
        n26525, n27101, n26524, n26523, n27100, n27099, n26770, 
        n26769, n26768, n26767, n26766, n26765, n26764, n26763, 
        n26762, n26761, n26760, n26759, n26758, n26757, n26756, 
        n26755, n26554, n26553, n26552;
    
    CCU2D sub_2078_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26550), .COUT(n26551));
    defparam sub_2078_add_2_25.INIT0 = 16'h5999;
    defparam sub_2078_add_2_25.INIT1 = 16'h5999;
    defparam sub_2078_add_2_25.INJECT1_0 = "NO";
    defparam sub_2078_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26549), .COUT(n26550));
    defparam sub_2078_add_2_23.INIT0 = 16'h5999;
    defparam sub_2078_add_2_23.INIT1 = 16'h5999;
    defparam sub_2078_add_2_23.INJECT1_0 = "NO";
    defparam sub_2078_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26548), .COUT(n26549));
    defparam sub_2078_add_2_21.INIT0 = 16'h5999;
    defparam sub_2078_add_2_21.INIT1 = 16'h5999;
    defparam sub_2078_add_2_21.INJECT1_0 = "NO";
    defparam sub_2078_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26547), .COUT(n26548));
    defparam sub_2078_add_2_19.INIT0 = 16'h5999;
    defparam sub_2078_add_2_19.INIT1 = 16'h5999;
    defparam sub_2078_add_2_19.INJECT1_0 = "NO";
    defparam sub_2078_add_2_19.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8332), .CK(debug_c_c), .CD(n31511), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2078_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26546), .COUT(n26547));
    defparam sub_2078_add_2_17.INIT0 = 16'h5999;
    defparam sub_2078_add_2_17.INIT1 = 16'h5999;
    defparam sub_2078_add_2_17.INJECT1_0 = "NO";
    defparam sub_2078_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26545), .COUT(n26546));
    defparam sub_2078_add_2_15.INIT0 = 16'h5999;
    defparam sub_2078_add_2_15.INIT1 = 16'h5999;
    defparam sub_2078_add_2_15.INJECT1_0 = "NO";
    defparam sub_2078_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26544), .COUT(n26545));
    defparam sub_2078_add_2_13.INIT0 = 16'h5999;
    defparam sub_2078_add_2_13.INIT1 = 16'h5999;
    defparam sub_2078_add_2_13.INJECT1_0 = "NO";
    defparam sub_2078_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26543), .COUT(n26544));
    defparam sub_2078_add_2_11.INIT0 = 16'h5999;
    defparam sub_2078_add_2_11.INIT1 = 16'h5999;
    defparam sub_2078_add_2_11.INJECT1_0 = "NO";
    defparam sub_2078_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26954), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_33.INIT1 = 16'h0000;
    defparam count_2676_add_4_33.INJECT1_0 = "NO";
    defparam count_2676_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26953), .COUT(n26954), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_31.INJECT1_0 = "NO";
    defparam count_2676_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26952), .COUT(n26953), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_29.INJECT1_0 = "NO";
    defparam count_2676_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26951), .COUT(n26952), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_27.INJECT1_0 = "NO";
    defparam count_2676_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26950), .COUT(n26951), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_25.INJECT1_0 = "NO";
    defparam count_2676_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26542), .COUT(n26543));
    defparam sub_2078_add_2_9.INIT0 = 16'h5999;
    defparam sub_2078_add_2_9.INIT1 = 16'h5999;
    defparam sub_2078_add_2_9.INJECT1_0 = "NO";
    defparam sub_2078_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26541), .COUT(n26542));
    defparam sub_2078_add_2_7.INIT0 = 16'h5999;
    defparam sub_2078_add_2_7.INIT1 = 16'h5999;
    defparam sub_2078_add_2_7.INJECT1_0 = "NO";
    defparam sub_2078_add_2_7.INJECT1_1 = "NO";
    FD1S3IX count_2676__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i0.GSR = "ENABLED";
    CCU2D count_2676_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26949), .COUT(n26950), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_23.INJECT1_0 = "NO";
    defparam count_2676_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26948), .COUT(n26949), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_21.INJECT1_0 = "NO";
    defparam count_2676_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26947), .COUT(n26948), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_19.INJECT1_0 = "NO";
    defparam count_2676_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26946), .COUT(n26947), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_17.INJECT1_0 = "NO";
    defparam count_2676_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26945), .COUT(n26946), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_15.INJECT1_0 = "NO";
    defparam count_2676_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26944), .COUT(n26945), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_13.INJECT1_0 = "NO";
    defparam count_2676_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26943), .COUT(n26944), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_11.INJECT1_0 = "NO";
    defparam count_2676_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26942), .COUT(n26943), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_9.INJECT1_0 = "NO";
    defparam count_2676_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26941), .COUT(n26942), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_7.INJECT1_0 = "NO";
    defparam count_2676_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26940), .COUT(n26941), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_5.INJECT1_0 = "NO";
    defparam count_2676_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26939), .COUT(n26940), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_3.INJECT1_0 = "NO";
    defparam count_2676_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27114), .S1(n8401));
    defparam sub_2081_add_2_33.INIT0 = 16'hf555;
    defparam sub_2081_add_2_33.INIT1 = 16'h0000;
    defparam sub_2081_add_2_33.INJECT1_0 = "NO";
    defparam sub_2081_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27113), .COUT(n27114));
    defparam sub_2081_add_2_31.INIT0 = 16'hf555;
    defparam sub_2081_add_2_31.INIT1 = 16'hf555;
    defparam sub_2081_add_2_31.INJECT1_0 = "NO";
    defparam sub_2081_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27112), .COUT(n27113));
    defparam sub_2081_add_2_29.INIT0 = 16'hf555;
    defparam sub_2081_add_2_29.INIT1 = 16'hf555;
    defparam sub_2081_add_2_29.INJECT1_0 = "NO";
    defparam sub_2081_add_2_29.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26939), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_1.INIT0 = 16'hF000;
    defparam count_2676_add_4_1.INIT1 = 16'h0555;
    defparam count_2676_add_4_1.INJECT1_0 = "NO";
    defparam count_2676_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27111), .COUT(n27112));
    defparam sub_2081_add_2_27.INIT0 = 16'hf555;
    defparam sub_2081_add_2_27.INIT1 = 16'hf555;
    defparam sub_2081_add_2_27.INJECT1_0 = "NO";
    defparam sub_2081_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27110), .COUT(n27111));
    defparam sub_2081_add_2_25.INIT0 = 16'hf555;
    defparam sub_2081_add_2_25.INIT1 = 16'hf555;
    defparam sub_2081_add_2_25.INJECT1_0 = "NO";
    defparam sub_2081_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27109), .COUT(n27110));
    defparam sub_2081_add_2_23.INIT0 = 16'hf555;
    defparam sub_2081_add_2_23.INIT1 = 16'hf555;
    defparam sub_2081_add_2_23.INJECT1_0 = "NO";
    defparam sub_2081_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27108), .COUT(n27109));
    defparam sub_2081_add_2_21.INIT0 = 16'hf555;
    defparam sub_2081_add_2_21.INIT1 = 16'hf555;
    defparam sub_2081_add_2_21.INJECT1_0 = "NO";
    defparam sub_2081_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27107), .COUT(n27108));
    defparam sub_2081_add_2_19.INIT0 = 16'hf555;
    defparam sub_2081_add_2_19.INIT1 = 16'hf555;
    defparam sub_2081_add_2_19.INJECT1_0 = "NO";
    defparam sub_2081_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27106), .COUT(n27107));
    defparam sub_2081_add_2_17.INIT0 = 16'hf555;
    defparam sub_2081_add_2_17.INIT1 = 16'hf555;
    defparam sub_2081_add_2_17.INJECT1_0 = "NO";
    defparam sub_2081_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27105), .COUT(n27106));
    defparam sub_2081_add_2_15.INIT0 = 16'hf555;
    defparam sub_2081_add_2_15.INIT1 = 16'hf555;
    defparam sub_2081_add_2_15.INJECT1_0 = "NO";
    defparam sub_2081_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26540), .COUT(n26541));
    defparam sub_2078_add_2_5.INIT0 = 16'h5999;
    defparam sub_2078_add_2_5.INIT1 = 16'h5999;
    defparam sub_2078_add_2_5.INJECT1_0 = "NO";
    defparam sub_2078_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27104), .COUT(n27105));
    defparam sub_2081_add_2_13.INIT0 = 16'hf555;
    defparam sub_2081_add_2_13.INIT1 = 16'hf555;
    defparam sub_2081_add_2_13.INJECT1_0 = "NO";
    defparam sub_2081_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26539), .COUT(n26540));
    defparam sub_2078_add_2_3.INIT0 = 16'h5999;
    defparam sub_2078_add_2_3.INIT1 = 16'h5999;
    defparam sub_2078_add_2_3.INJECT1_0 = "NO";
    defparam sub_2078_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26539));
    defparam sub_2078_add_2_1.INIT0 = 16'h0000;
    defparam sub_2078_add_2_1.INIT1 = 16'h5999;
    defparam sub_2078_add_2_1.INJECT1_0 = "NO";
    defparam sub_2078_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26538), .S1(n8367));
    defparam sub_2080_add_2_33.INIT0 = 16'h5999;
    defparam sub_2080_add_2_33.INIT1 = 16'h0000;
    defparam sub_2080_add_2_33.INJECT1_0 = "NO";
    defparam sub_2080_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26537), .COUT(n26538));
    defparam sub_2080_add_2_31.INIT0 = 16'h5999;
    defparam sub_2080_add_2_31.INIT1 = 16'h5999;
    defparam sub_2080_add_2_31.INJECT1_0 = "NO";
    defparam sub_2080_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26536), .COUT(n26537));
    defparam sub_2080_add_2_29.INIT0 = 16'h5999;
    defparam sub_2080_add_2_29.INIT1 = 16'h5999;
    defparam sub_2080_add_2_29.INJECT1_0 = "NO";
    defparam sub_2080_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26535), .COUT(n26536));
    defparam sub_2080_add_2_27.INIT0 = 16'h5999;
    defparam sub_2080_add_2_27.INIT1 = 16'h5999;
    defparam sub_2080_add_2_27.INJECT1_0 = "NO";
    defparam sub_2080_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26534), .COUT(n26535));
    defparam sub_2080_add_2_25.INIT0 = 16'h5999;
    defparam sub_2080_add_2_25.INIT1 = 16'h5999;
    defparam sub_2080_add_2_25.INJECT1_0 = "NO";
    defparam sub_2080_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27103), .COUT(n27104));
    defparam sub_2081_add_2_11.INIT0 = 16'hf555;
    defparam sub_2081_add_2_11.INIT1 = 16'hf555;
    defparam sub_2081_add_2_11.INJECT1_0 = "NO";
    defparam sub_2081_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26533), .COUT(n26534));
    defparam sub_2080_add_2_23.INIT0 = 16'h5999;
    defparam sub_2080_add_2_23.INIT1 = 16'h5999;
    defparam sub_2080_add_2_23.INJECT1_0 = "NO";
    defparam sub_2080_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26532), .COUT(n26533));
    defparam sub_2080_add_2_21.INIT0 = 16'h5999;
    defparam sub_2080_add_2_21.INIT1 = 16'h5999;
    defparam sub_2080_add_2_21.INJECT1_0 = "NO";
    defparam sub_2080_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27102), .COUT(n27103));
    defparam sub_2081_add_2_9.INIT0 = 16'hf555;
    defparam sub_2081_add_2_9.INIT1 = 16'hf555;
    defparam sub_2081_add_2_9.INJECT1_0 = "NO";
    defparam sub_2081_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26531), .COUT(n26532));
    defparam sub_2080_add_2_19.INIT0 = 16'h5999;
    defparam sub_2080_add_2_19.INIT1 = 16'h5999;
    defparam sub_2080_add_2_19.INJECT1_0 = "NO";
    defparam sub_2080_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26530), .COUT(n26531));
    defparam sub_2080_add_2_17.INIT0 = 16'h5999;
    defparam sub_2080_add_2_17.INIT1 = 16'h5999;
    defparam sub_2080_add_2_17.INJECT1_0 = "NO";
    defparam sub_2080_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26529), .COUT(n26530));
    defparam sub_2080_add_2_15.INIT0 = 16'h5999;
    defparam sub_2080_add_2_15.INIT1 = 16'h5999;
    defparam sub_2080_add_2_15.INJECT1_0 = "NO";
    defparam sub_2080_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26528), .COUT(n26529));
    defparam sub_2080_add_2_13.INIT0 = 16'h5999;
    defparam sub_2080_add_2_13.INIT1 = 16'h5999;
    defparam sub_2080_add_2_13.INJECT1_0 = "NO";
    defparam sub_2080_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26527), .COUT(n26528));
    defparam sub_2080_add_2_11.INIT0 = 16'h5999;
    defparam sub_2080_add_2_11.INIT1 = 16'h5999;
    defparam sub_2080_add_2_11.INJECT1_0 = "NO";
    defparam sub_2080_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26526), .COUT(n26527));
    defparam sub_2080_add_2_9.INIT0 = 16'h5999;
    defparam sub_2080_add_2_9.INIT1 = 16'h5999;
    defparam sub_2080_add_2_9.INJECT1_0 = "NO";
    defparam sub_2080_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26525), .COUT(n26526));
    defparam sub_2080_add_2_7.INIT0 = 16'h5999;
    defparam sub_2080_add_2_7.INIT1 = 16'h5999;
    defparam sub_2080_add_2_7.INJECT1_0 = "NO";
    defparam sub_2080_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27101), .COUT(n27102));
    defparam sub_2081_add_2_7.INIT0 = 16'hf555;
    defparam sub_2081_add_2_7.INIT1 = 16'hf555;
    defparam sub_2081_add_2_7.INJECT1_0 = "NO";
    defparam sub_2081_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2080_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26524), .COUT(n26525));
    defparam sub_2080_add_2_5.INIT0 = 16'h5999;
    defparam sub_2080_add_2_5.INIT1 = 16'h5999;
    defparam sub_2080_add_2_5.INJECT1_0 = "NO";
    defparam sub_2080_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26523), .COUT(n26524));
    defparam sub_2080_add_2_3.INIT0 = 16'h5999;
    defparam sub_2080_add_2_3.INIT1 = 16'h5999;
    defparam sub_2080_add_2_3.INJECT1_0 = "NO";
    defparam sub_2080_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2080_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26523));
    defparam sub_2080_add_2_1.INIT0 = 16'h0000;
    defparam sub_2080_add_2_1.INIT1 = 16'h5999;
    defparam sub_2080_add_2_1.INJECT1_0 = "NO";
    defparam sub_2080_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27100), .COUT(n27101));
    defparam sub_2081_add_2_5.INIT0 = 16'hf555;
    defparam sub_2081_add_2_5.INIT1 = 16'hf555;
    defparam sub_2081_add_2_5.INJECT1_0 = "NO";
    defparam sub_2081_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27099), .COUT(n27100));
    defparam sub_2081_add_2_3.INIT0 = 16'hf555;
    defparam sub_2081_add_2_3.INIT1 = 16'hf555;
    defparam sub_2081_add_2_3.INJECT1_0 = "NO";
    defparam sub_2081_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27099));
    defparam sub_2081_add_2_1.INIT0 = 16'h0000;
    defparam sub_2081_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2081_add_2_1.INJECT1_0 = "NO";
    defparam sub_2081_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31409), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31409), .PD(n16842), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26770), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26769), .COUT(n26770), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26768), .COUT(n26769), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26767), .COUT(n26768), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26766), .COUT(n26767), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26765), .COUT(n26766), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26764), .COUT(n26765), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26763), .COUT(n26764), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26762), .COUT(n26763), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26761), .COUT(n26762), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26760), .COUT(n26761), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26759), .COUT(n26760), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26758), .COUT(n26759), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26757), .COUT(n26758), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26756), .COUT(n26757), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26755), .COUT(n26756), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26755), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1S3IX count_2676__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i1.GSR = "ENABLED";
    FD1S3IX count_2676__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i2.GSR = "ENABLED";
    FD1S3IX count_2676__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i3.GSR = "ENABLED";
    FD1S3IX count_2676__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i4.GSR = "ENABLED";
    FD1S3IX count_2676__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i5.GSR = "ENABLED";
    FD1S3IX count_2676__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i6.GSR = "ENABLED";
    FD1S3IX count_2676__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i7.GSR = "ENABLED";
    FD1S3IX count_2676__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i8.GSR = "ENABLED";
    FD1S3IX count_2676__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i9.GSR = "ENABLED";
    FD1S3IX count_2676__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i10.GSR = "ENABLED";
    FD1S3IX count_2676__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i11.GSR = "ENABLED";
    FD1S3IX count_2676__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i12.GSR = "ENABLED";
    FD1S3IX count_2676__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i13.GSR = "ENABLED";
    FD1S3IX count_2676__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i14.GSR = "ENABLED";
    FD1S3IX count_2676__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i15.GSR = "ENABLED";
    FD1S3IX count_2676__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i16.GSR = "ENABLED";
    FD1S3IX count_2676__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i17.GSR = "ENABLED";
    FD1S3IX count_2676__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i18.GSR = "ENABLED";
    FD1S3IX count_2676__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i19.GSR = "ENABLED";
    FD1S3IX count_2676__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i20.GSR = "ENABLED";
    FD1S3IX count_2676__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i21.GSR = "ENABLED";
    FD1S3IX count_2676__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i22.GSR = "ENABLED";
    FD1S3IX count_2676__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i23.GSR = "ENABLED";
    FD1S3IX count_2676__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i24.GSR = "ENABLED";
    FD1S3IX count_2676__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i25.GSR = "ENABLED";
    FD1S3IX count_2676__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i26.GSR = "ENABLED";
    FD1S3IX count_2676__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i27.GSR = "ENABLED";
    FD1S3IX count_2676__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i28.GSR = "ENABLED";
    FD1S3IX count_2676__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i29.GSR = "ENABLED";
    FD1S3IX count_2676__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i30.GSR = "ENABLED";
    FD1S3IX count_2676__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i31.GSR = "ENABLED";
    CCU2D sub_2078_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26554), .S1(n8332));
    defparam sub_2078_add_2_33.INIT0 = 16'h5555;
    defparam sub_2078_add_2_33.INIT1 = 16'h0000;
    defparam sub_2078_add_2_33.INJECT1_0 = "NO";
    defparam sub_2078_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26553), .COUT(n26554));
    defparam sub_2078_add_2_31.INIT0 = 16'h5999;
    defparam sub_2078_add_2_31.INIT1 = 16'h5999;
    defparam sub_2078_add_2_31.INJECT1_0 = "NO";
    defparam sub_2078_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26552), .COUT(n26553));
    defparam sub_2078_add_2_29.INIT0 = 16'h5999;
    defparam sub_2078_add_2_29.INIT1 = 16'h5999;
    defparam sub_2078_add_2_29.INJECT1_0 = "NO";
    defparam sub_2078_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2078_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26551), .COUT(n26552));
    defparam sub_2078_add_2_27.INIT0 = 16'h5999;
    defparam sub_2078_add_2_27.INIT1 = 16'h5999;
    defparam sub_2078_add_2_27.INJECT1_0 = "NO";
    defparam sub_2078_add_2_27.INJECT1_1 = "NO";
    
endmodule
