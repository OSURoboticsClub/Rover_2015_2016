// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Thu Apr  7 06:49:37 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    output expansion4 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire n32376 /* synthesis nomerge= */ ;
    
    wire GND_net, VCC_net, uart_rx_c, n10643, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, signal_light_c, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
        encoder_la_c, encoder_lb_c, encoder_li_c, rc_ch1_c, rc_ch2_c, 
        rc_ch3_c, rc_ch4_c, rc_ch7_c, rc_ch8_c, motor_pwm_l_c, xbee_pause_c, 
        debug_c_7, debug_c_5, debug_c_4, debug_c_3, debug_c_2, debug_c_0;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire rw, n14121, n14013, n13918;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    
    wire n17, n6, n26485, n24, n26592, n13269, n34, n28853, 
        n26486;
    wire [7:0]n8262;
    
    wire n26604, n22;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n12, n20681, n20679, n14, n20671, n20670, n13;
    wire [31:0]n1295;
    
    wire n26607, n22_adj_523, n28765, n28775, n5632, n8129, n2673, 
        n3892, n13624, n8, n9118;
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[12:21])
    
    wire n46, n27462, n28770, n3, n30331, n5, n3_adj_524, n28421, 
        n17_adj_525;
    wire [2:0]read_size_adj_852;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(93[12:21])
    
    wire n28723, n13594, n13589;
    wire [15:0]n281;
    
    wire n6_adj_527, n30330, n32, n32_adj_528, n13574, n241;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire step_clk, prev_step_clk;
    wire [31:0]read_value_adj_858;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_859;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select, n6_adj_563, n2644, n302, n13534;
    wire [31:0]n580;
    
    wire n1;
    wire [7:0]control_reg_adj_867;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_868;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_869;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire fault_latched, step_clk_adj_565, prev_step_clk_adj_566;
    wire [31:0]read_value_adj_870;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_871;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_601, n28910, n28148, n3_adj_602, n6_adj_603, 
        n19;
    wire [31:0]n580_adj_890;
    
    wire n16;
    wire [7:0]control_reg_adj_908;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_909;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_910;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire int_step, step_clk_adj_605, prev_step_clk_adj_606;
    wire [31:0]read_value_adj_911;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_912;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_641, n12_adj_642;
    wire [31:0]n99_adj_1268;
    
    wire n28017, n28137;
    wire [7:0]n571_adj_930;
    
    wire n19585;
    wire [7:0]control_reg_adj_949;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_951;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping;
    wire [31:0]read_value_adj_952;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_953;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_678, n28172, n19_adj_679, n3_adj_680, n8_adj_681;
    wire [31:0]n99_adj_1273;
    
    wire n16_adj_682, n12_adj_683, n11, n32377, n20668;
    wire [3:0]n32520;
    
    wire n28748, qreset;
    wire [31:0]read_value_adj_993;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[13:23])
    wire [2:0]read_size_adj_994;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(67[12:21])
    
    wire prev_select_adj_719, n47, n21563, n21310;
    wire [31:0]\register[1]_adj_1000 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    wire [31:0]read_value_adj_1002;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[13:23])
    wire [2:0]read_size_adj_1003;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(67[12:21])
    
    wire prev_select_adj_754, n176, n28670, n28196, n6_adj_755, n3806, 
        n6_adj_756, n6_adj_757, n8_adj_758, n5_adj_759, n2, n4, 
        n2_adj_760, n1_adj_761, n8_adj_762, n5_adj_763, n2_adj_764, 
        n2_adj_765, n5_adj_766;
    wire [14:0]n66_adj_1398;
    
    wire n8_adj_767, n2_adj_768, n5_adj_769, n2_adj_770, n5_adj_771, 
        n8_adj_772, n5_adj_773, n8_adj_774, n2_adj_775, n5_adj_776, 
        n8_adj_777, n3_adj_778, n3_adj_779, n30324, n6_adj_780, n6_adj_781, 
        n3_adj_782, n3_adj_783, n6_adj_784, n6_adj_785, n3_adj_786, 
        n6_adj_787, n3_adj_788, n6_adj_789, n3_adj_790, n6_adj_791, 
        n3_adj_792, n6_adj_793, n3_adj_794, n6_adj_795, n6_adj_796, 
        n6_adj_797, n3_adj_798, n6_adj_799, n3_adj_800, n3_adj_801, 
        n3_adj_802, n6_adj_803, n3_adj_804, n6_adj_805, n6_adj_806, 
        n3_adj_807, n6_adj_808, n21533, n30321, n30317, n3_adj_809, 
        n6_adj_810, n30316, n30314, n30313, n30311, n30310, n30307, 
        n3_adj_811, n6_adj_812, n25973, n25972, n28851, n25971, 
        n3_adj_813, n30491, n30489, n30488, n14309, n14308, n14307, 
        n14306;
    wire [31:0]n6891;
    
    wire n13_adj_814, n25970, n30479, n30478;
    wire [7:0]n8271;
    
    wire n25969, n25968, n25967, n11_adj_815, n11_adj_816, n28218, 
        n14291, n26618, n30305, n22_adj_817, n30, n14284, n6_adj_818;
    wire [3:0]state_adj_1038;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    
    wire select_clk, n30463, n8894, n28672, n30454, n8890, n30445, 
        n30444, n28671, n26601, n4_adj_819, n30427, n30422, n30421, 
        n28857, n30417, n30413, n4_adj_820, n20944, n4_adj_821, 
        n30411, n3989, n3666, n26465, n32386, n3_adj_822;
    wire [2:0]quadA_delayed_adj_1102;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [2:0]quadB_delayed_adj_1103;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n30406, n26787, n3_adj_823, n28323, n28725, n26671, n9136, 
        n9128, n32385, n9125, n9122, n28859, n32384, n30398, n30396, 
        n30395, n30394, n30391, n2_adj_826, n30385, n31, n19_adj_827, 
        n30383, n32383, n30380, n30379, n30303, n32382, n26596, 
        n26484, n28605, n32381, n30374, n30373, n30372, n30371, 
        n30370, n30367, n30366, n28324, n30361, n7504, n32380, 
        n28184, n30358, n30350, n30349, n26299, n32379, n30344, 
        n28522, n30342, n30340, n30339, n107, n28855, n26585, 
        n30338, n28773, n26507;
    
    VHI i2 (.Z(VCC_net));
    GlobalControlPeripheral global_control (.debug_c_c(debug_c_c), .n32384(n32384), 
            .\databus[1] (databus[1]), .\select[1] (select[1]), .rw(rw), 
            .n46(n46), .n32381(n32381), .read_size({read_size}), .n30307(n30307), 
            .n302(n302), .n26507(n26507), .n30330(n30330), .n32380(n32380), 
            .n32385(n32385), .\register_addr[4] (register_addr[4]), .\register_addr[3] (register_addr[3]), 
            .n21310(n21310), .xbee_pause_c(xbee_pause_c), .\register_addr[0] (register_addr[0]), 
            .n9118(n9118), .n30478(n30478), .n11(n11_adj_816), .\register_addr[1] (register_addr[1]), 
            .n30366(n30366), .n30413(n30413), .\register_addr[2] (register_addr[2]), 
            .n6(n6_adj_527), .n30491(n30491), .n28421(n28421), .n30395(n30395), 
            .n176(n176), .n8(n8_adj_681), .\control_reg[7] (control_reg_adj_908[7]), 
            .n26486(n26486), .n32(n32_adj_528), .\control_reg[7]_adj_228 (control_reg_adj_867[7]), 
            .n26485(n26485), .n32_adj_229(n32), .\control_reg[7]_adj_230 (control_reg_adj_949[7]), 
            .n26585(n26585), .stepping(stepping), .\control_reg[7]_adj_231 (control_reg[7]), 
            .n26484(n26484), .n34(n34), .\state[0] (state_adj_1038[0]), 
            .n22(n22_adj_817), .n27462(n27462), .signal_light_c(signal_light_c), 
            .n31(n31), .n19(n19_adj_827), .n28218(n28218), .n30344(n30344), 
            .n30417(n30417), .n13594(n13594), .n32377(n32377), .\select[3] (select[3]), 
            .n30358(n30358), .\register_addr[5] (register_addr[5]), .n30361(n30361), 
            .read_value({read_value}), .GND_net(GND_net), .n30394(n30394), 
            .n30324(n30324), .n30489(n30489), .n8890(n8890)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(495[45] 505[74])
    LUT4 i14569_2_lut (.A(reset_count[11]), .B(reset_count[13]), .Z(n20944)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i14569_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_307_3_lut_4_lut (.A(n30398), .B(register_addr[5]), 
         .C(n32379), .D(prev_select_adj_601), .Z(n30316)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i1_2_lut_rep_307_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(n30398), .B(register_addr[5]), .C(n32380), 
         .D(prev_select_adj_601), .Z(n14121)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 Select_4204_i3_2_lut_3_lut_4_lut (.A(n30398), .B(register_addr[5]), 
         .C(read_value_adj_870[13]), .D(rw), .Z(n3_adj_783)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4204_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i14892_2_lut_2_lut (.A(n32380), .B(databus[2]), .Z(n580_adj_890[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14892_2_lut_2_lut.init = 16'h4444;
    LUT4 Select_4210_i3_2_lut_3_lut_4_lut (.A(n30398), .B(register_addr[5]), 
         .C(read_value_adj_870[11]), .D(rw), .Z(n3_adj_782)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4210_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4213_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[10]), 
         .D(n32379), .Z(n3_adj_778)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4213_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4216_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[9]), 
         .D(n32379), .Z(n3_adj_788)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4216_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4150_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[31]), 
         .D(n32379), .Z(n3_adj_823)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4150_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4153_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[30]), 
         .D(rw), .Z(n3_adj_822)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4153_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4156_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[29]), 
         .D(rw), .Z(n3_adj_524)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4156_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4159_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[28]), 
         .D(rw), .Z(n3_adj_602)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4159_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4162_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[27]), 
         .D(rw), .Z(n3_adj_809)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4162_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4165_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[26]), 
         .D(rw), .Z(n3_adj_680)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4165_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4168_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[25]), 
         .D(rw), .Z(n3_adj_811)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4168_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4171_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[24]), 
         .D(rw), .Z(n3_adj_807)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4171_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i21519 (.BLUT(n28670), .ALUT(n28671), .C0(register_addr[0]), 
          .Z(n28672));
    LUT4 Select_4174_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[23]), 
         .D(rw), .Z(n3_adj_813)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4174_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_4_lut (.A(register_addr[1]), .B(div_factor_reg_adj_868[20]), 
         .C(steps_reg_adj_869[20]), .D(register_addr[0]), .Z(n12_adj_642)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 Select_4177_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[22]), 
         .D(rw), .Z(n3_adj_800)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4177_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4180_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[21]), 
         .D(rw), .Z(n3)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4180_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4183_i3_2_lut_3_lut_4_lut (.A(n30398), .B(register_addr[5]), 
         .C(read_value_adj_870[20]), .D(rw), .Z(n3_adj_801)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4183_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4186_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[19]), 
         .D(rw), .Z(n3_adj_798)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4186_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4189_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[18]), 
         .D(rw), .Z(n3_adj_794)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4189_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4192_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[17]), 
         .D(rw), .Z(n3_adj_804)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4192_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4195_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[16]), 
         .D(rw), .Z(n3_adj_802)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4195_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4198_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[15]), 
         .D(rw), .Z(n3_adj_792)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4198_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4201_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[14]), 
         .D(rw), .Z(n3_adj_790)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4201_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4207_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[12]), 
         .D(rw), .Z(n3_adj_779)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4207_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4219_i3_2_lut_3_lut_4_lut (.A(n30398), .B(n32377), .C(read_value_adj_870[8]), 
         .D(rw), .Z(n3_adj_786)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam Select_4219_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i15_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n30413), .C(rw), 
         .D(select[3]), .Z(n47)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam i15_2_lut_3_lut_4_lut.init = 16'hd000;
    LUT4 i114_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n30413), .C(prev_select_adj_719), 
         .D(select[3]), .Z(n14291)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam i114_2_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i15_2_lut_rep_330_3_lut_4_lut (.A(register_addr[4]), .B(n30413), 
         .C(n32379), .D(select[3]), .Z(n30339)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam i15_2_lut_rep_330_3_lut_4_lut.init = 16'h2000;
    LUT4 i114_2_lut_3_lut_4_lut_adj_458 (.A(register_addr[4]), .B(n30413), 
         .C(prev_select_adj_754), .D(select[3]), .Z(n13589)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam i114_2_lut_3_lut_4_lut_adj_458.init = 16'h0200;
    LUT4 i1_2_lut_rep_296_3_lut_3_lut (.A(n32380), .B(select_clk), .C(n8129), 
         .Z(n30305)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_296_3_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_435 (.A(reset_count[7]), .B(reset_count[8]), .Z(n30444)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i1_2_lut_rep_435.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(reset_count[7]), .B(reset_count[8]), .C(reset_count[6]), 
         .D(reset_count[5]), .Z(n4_adj_819)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i1_3_lut_4_lut.init = 16'hfe00;
    LUT4 i21853_4_lut_rep_486 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n32380)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_486.init = 16'h23af;
    LUT4 Select_4225_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[2]), 
         .D(rw), .Z(n2)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4225_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4222_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[5]), 
         .D(rw), .Z(n2_adj_768)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4222_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4220_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[7]), 
         .D(rw), .Z(n2_adj_775)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4220_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i21853_4_lut_rep_487 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n32381)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_487.init = 16'h23af;
    LUT4 Select_4223_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[4]), 
         .D(n32379), .Z(n2_adj_826)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4223_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4221_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[6]), 
         .D(rw), .Z(n2_adj_770)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4221_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4224_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[3]), 
         .D(rw), .Z(n2_adj_765)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4224_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4226_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[1]), 
         .D(rw), .Z(n2_adj_760)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4226_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4227_i2_2_lut_3_lut_4_lut (.A(n30427), .B(n30479), .C(read_value_adj_911[0]), 
         .D(rw), .Z(n2_adj_764)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4227_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_adj_459 (.A(n30427), .B(n30479), .C(n32380), 
         .D(prev_select_adj_641), .Z(n13918)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_adj_459.init = 16'h0002;
    LUT4 i1_2_lut_rep_335_3_lut_4_lut (.A(n30427), .B(n30479), .C(n32379), 
         .D(prev_select_adj_641), .Z(n30344)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_rep_335_3_lut_4_lut.init = 16'h0002;
    LUT4 i21853_4_lut_rep_488 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n32382)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_488.init = 16'h23af;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_adj_460 (.A(n30427), .B(n30488), .C(n32380), 
         .D(prev_select), .Z(n2644)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_adj_460.init = 16'h0002;
    LUT4 i1_2_lut_rep_315_3_lut_4_lut (.A(n30427), .B(n30488), .C(n32379), 
         .D(prev_select), .Z(n30324)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_rep_315_3_lut_4_lut.init = 16'h0002;
    LUT4 Select_4226_i4_2_lut_3_lut_4_lut (.A(n30427), .B(n30488), .C(read_value_adj_858[1]), 
         .D(rw), .Z(n4)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4226_i4_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i21853_4_lut_rep_489 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n32383)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_489.init = 16'h23af;
    LUT4 i173_2_lut_rep_454 (.A(reset_count[10]), .B(reset_count[9]), .Z(n30463)) /* synthesis lut_function=(A (B)) */ ;
    defparam i173_2_lut_rep_454.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_461 (.A(reset_count[10]), .B(reset_count[9]), 
         .C(reset_count[14]), .D(reset_count[4]), .Z(n26465)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_461.init = 16'h8000;
    LUT4 i21853_4_lut_rep_490 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n32384)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_490.init = 16'h23af;
    FD1P3AX reset_count_2606_2607__i1 (.D(n66_adj_1398[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i1.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_4_lut_3_lut_4_lut (.A(n32380), .B(state_adj_1038[0]), 
         .C(n8129), .D(select_clk), .Z(n32520[0])) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hcc9c;
    LUT4 i21853_4_lut_rep_491 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n32385)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_491.init = 16'h23af;
    LUT4 i1_2_lut_rep_470 (.A(register_addr[4]), .B(n32377), .Z(n30479)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i1_2_lut_rep_470.init = 16'hbbbb;
    LUT4 i21452_4_lut (.A(n28522), .B(n20944), .C(n30463), .D(n30444), 
         .Z(n28605)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i21452_4_lut.init = 16'hfcec;
    LUT4 i21374_3_lut (.A(reset_count[5]), .B(reset_count[6]), .C(reset_count[4]), 
         .Z(n28522)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i21374_3_lut.init = 16'hc8c8;
    LUT4 i1_2_lut_rep_358_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(rw), .D(n30427), .Z(n30367)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i1_2_lut_rep_358_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_2_lut_rep_364_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(prev_select_adj_641), .D(n30427), .Z(n30373)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i2_2_lut_rep_364_3_lut_4_lut.init = 16'h0400;
    LUT4 i21853_4_lut_rep_492 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n32386)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_492.init = 16'h23af;
    LUT4 i2_4_lut_4_lut (.A(n32380), .B(n28184), .C(n30491), .D(n30338), 
         .Z(n9136)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (D)))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h5100;
    LUT4 i1_4_lut_adj_462 (.A(div_factor_reg_adj_909[9]), .B(register_addr[1]), 
         .C(steps_reg_adj_910[9]), .D(register_addr[0]), .Z(n28148)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_462.init = 16'hc088;
    LUT4 i21645_2_lut (.A(int_step), .B(control_reg_adj_908[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i21645_2_lut.init = 16'h9999;
    LUT4 i14565_2_lut_2_lut (.A(n32380), .B(databus[4]), .Z(n580[4])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14565_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_479 (.A(register_addr[4]), .B(n32377), .Z(n30488)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i1_2_lut_rep_479.init = 16'heeee;
    LUT4 i1_2_lut_rep_363_3_lut_4_lut (.A(register_addr[4]), .B(n32377), 
         .C(rw), .D(n30427), .Z(n30372)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i1_2_lut_rep_363_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_2_lut_3_lut (.A(register_addr[4]), .B(register_addr[5]), .C(register_addr[3]), 
         .Z(n6_adj_527)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i2_2_lut_3_lut.init = 16'hfefe;
    LUT4 i2_2_lut_rep_341_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(prev_select), .D(n30427), .Z(n30350)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i2_2_lut_rep_341_3_lut_4_lut.init = 16'h0100;
    LUT4 Select_4195_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[16]), 
         .D(rw), .Z(n6_adj_803)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4195_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_2_lut (.A(n32380), .B(n8129), .Z(n107)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 Select_4198_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[15]), 
         .D(rw), .Z(n6_adj_793)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4198_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i3_4_lut (.A(n30316), .B(n28196), .C(register_addr[5]), .D(n30411), 
         .Z(n8894)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(526[4] 555[11])
    defparam i3_4_lut.init = 16'h0800;
    LUT4 i2_4_lut_4_lut_adj_463 (.A(n32380), .B(n28196), .C(n30413), .D(n30331), 
         .Z(n9128)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (D)))) */ ;
    defparam i2_4_lut_4_lut_adj_463.init = 16'h5100;
    LUT4 Select_4201_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[14]), 
         .D(n32379), .Z(n6_adj_791)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4201_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i15130_2_lut_2_lut (.A(n32380), .B(databus[0]), .Z(n571_adj_930[0])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15130_2_lut_2_lut.init = 16'h4444;
    LUT4 i14515_2_lut_2_lut (.A(n32380), .B(n7504), .Z(n241)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14515_2_lut_2_lut.init = 16'h4444;
    PFUMX i14297 (.BLUT(n20671), .ALUT(n13), .C0(register_addr[0]), .Z(n6891[6]));
    LUT4 i29_4_lut (.A(n28017), .B(reset_count[14]), .C(n30444), .D(n30463), 
         .Z(n16)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i29_4_lut.init = 16'hca0a;
    LUT4 i2_4_lut (.A(n20944), .B(n30463), .C(reset_count[12]), .D(n4_adj_819), 
         .Z(n19)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i2_4_lut.init = 16'hfefa;
    PFUMX i14294 (.BLUT(n20668), .ALUT(n12), .C0(register_addr[0]), .Z(n20670));
    LUT4 i2_4_lut_adj_464 (.A(n20944), .B(reset_count[12]), .C(n26465), 
         .D(reset_count[6]), .Z(n28017)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i2_4_lut_adj_464.init = 16'h1000;
    LUT4 Select_4207_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[12]), 
         .D(n32379), .Z(n6_adj_781)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4207_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21853_4_lut_rep_333 (.A(reset_count[5]), .B(reset_count[14]), 
         .C(n16), .D(n19), .Z(n30342)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i21853_4_lut_rep_333.init = 16'h23af;
    LUT4 Select_4219_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[8]), 
         .D(n32379), .Z(n6_adj_787)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4219_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21517_3_lut (.A(Stepper_Y_M1_c_1), .B(div_factor_reg_adj_868[1]), 
         .C(register_addr[1]), .Z(n28670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21517_3_lut.init = 16'hcaca;
    LUT4 Select_4227_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[0]), 
         .D(n32379), .Z(n8_adj_762)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4227_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21518_3_lut (.A(fault_latched), .B(steps_reg_adj_869[1]), .C(register_addr[1]), 
         .Z(n28671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21518_3_lut.init = 16'hcaca;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB encoder_li_pad (.I(encoder_li), .O(encoder_li_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    IB encoder_lb_pad (.I(encoder_lb), .O(encoder_lb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    IB encoder_la_pad (.I(encoder_la), .O(encoder_la_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    IB encoder_ri_pad (.I(encoder_ri), .O(encoder_ri_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    IB encoder_rb_pad (.I(encoder_rb), .O(encoder_rb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    IB encoder_ra_pad (.I(encoder_ra), .O(encoder_ra_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    IB uart_rx_pad (.I(uart_rx), .O(uart_rx_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    OB debug_pad_0 (.I(debug_c_0), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_1 (.I(n10643), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_6 (.I(n32380), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB motor_pwm_r_pad (.I(GND_net), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    OB expansion5_pad (.I(GND_net), .O(expansion5));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    OB expansion4_pad (.I(GND_net), .O(expansion4));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    OB expansion3_pad (.I(GND_net), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    OB expansion2_pad (.I(GND_net), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion1_pad (.I(GND_net), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB uart_tx_pad (.I(n10643), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    CCU2D reset_count_2606_2607_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25973), .S0(n66_adj_1398[13]), 
          .S1(n66_adj_1398[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2606_2607_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25972), .COUT(n25973), .S0(n66_adj_1398[11]), 
          .S1(n66_adj_1398[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2606_2607_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25971), .COUT(n25972), .S0(n66_adj_1398[9]), 
          .S1(n66_adj_1398[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2606_2607_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25970), .COUT(n25971), .S0(n66_adj_1398[7]), 
          .S1(n66_adj_1398[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2606_2607_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25969), .COUT(n25970), .S0(n66_adj_1398[5]), 
          .S1(n66_adj_1398[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_7.INJECT1_1 = "NO";
    CCU2D reset_count_2606_2607_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25968), .COUT(n25969), .S0(n66_adj_1398[3]), 
          .S1(n66_adj_1398[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_5.INJECT1_1 = "NO";
    LUT4 i2_3_lut_3_lut_4_lut (.A(prev_select), .B(n30396), .C(n11_adj_816), 
         .D(n32380), .Z(n9125)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_3_lut_3_lut_4_lut.init = 16'h0040;
    CCU2D reset_count_2606_2607_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25967), .COUT(n25968), .S0(n66_adj_1398[1]), 
          .S1(n66_adj_1398[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2606_2607_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2606_2607_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n25967), .S1(n66_adj_1398[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2606_2607_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2606_2607_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2606_2607_add_4_1.INJECT1_1 = "NO";
    LUT4 i14872_2_lut_2_lut (.A(n32380), .B(databus[7]), .Z(n281[15])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14872_2_lut_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_3_lut (.A(n30383), .B(n1295[17]), .C(n1295[20]), .Z(n26671)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i2_3_lut_3_lut.init = 16'hfdfd;
    FD1P3AX reset_count_2606_2607__i2 (.D(n66_adj_1398[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i2.GSR = "ENABLED";
    LUT4 i21688_4_lut_4_lut (.A(n30383), .B(n4_adj_821), .C(n5632), .D(n1295[14]), 
         .Z(n13574)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i21688_4_lut_4_lut.init = 16'h2a00;
    LUT4 i3_4_lut_adj_465 (.A(n26299), .B(n30463), .C(reset_count[11]), 
         .D(reset_count[8]), .Z(n26787)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_465.init = 16'hc080;
    LUT4 i2_3_lut (.A(reset_count[5]), .B(reset_count[7]), .C(reset_count[6]), 
         .Z(n26299)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_rep_331_4_lut (.A(select[3]), .B(n30385), .C(n30379), 
         .D(prev_select_adj_719), .Z(n30340)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam i2_3_lut_rep_331_4_lut.init = 16'h0020;
    LUT4 Select_4210_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[11]), 
         .D(rw), .Z(n6_adj_784)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4210_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4204_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[13]), 
         .D(rw), .Z(n6_adj_785)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4204_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_rep_312_4_lut (.A(select[3]), .B(n30385), .C(n30406), 
         .D(prev_select_adj_754), .Z(n30321)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam i2_3_lut_rep_312_4_lut.init = 16'h0080;
    LUT4 i105_4_lut (.A(n11), .B(sendcount[0]), .C(n16_adj_682), .D(n12_adj_683), 
         .Z(n17_adj_525)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    defparam i105_4_lut.init = 16'h3336;
    LUT4 i1_4_lut_adj_466 (.A(n19585), .B(div_factor_reg_adj_868[24]), .C(steps_reg_adj_869[24]), 
         .D(register_addr[0]), .Z(n99_adj_1273[24])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_466.init = 16'ha088;
    GSR GSR_INST (.GSR(VCC_net));
    FD1P3AX reset_count_2606_2607__i3 (.D(n66_adj_1398[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i4 (.D(n66_adj_1398[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i5 (.D(n66_adj_1398[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i6 (.D(n66_adj_1398[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i7 (.D(n66_adj_1398[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i8 (.D(n66_adj_1398[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i9 (.D(n66_adj_1398[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i10 (.D(n66_adj_1398[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i11 (.D(n66_adj_1398[10]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i12 (.D(n66_adj_1398[11]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i13 (.D(n66_adj_1398[12]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i14 (.D(n66_adj_1398[13]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2606_2607__i15 (.D(n66_adj_1398[14]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2606_2607__i15.GSR = "ENABLED";
    LUT4 Select_4213_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[10]), 
         .D(rw), .Z(n6_adj_780)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4213_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4216_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[9]), 
         .D(rw), .Z(n6_adj_789)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4216_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4220_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[7]), 
         .D(rw), .Z(n8_adj_777)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4220_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4221_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[6]), 
         .D(n32379), .Z(n8_adj_774)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4221_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4222_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[5]), 
         .D(rw), .Z(n8_adj_767)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4222_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4223_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[4]), 
         .D(rw), .Z(n8_adj_772)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4223_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    VLO i1 (.Z(GND_net));
    EncoderPeripheral_U11 left_encoder (.prev_select(prev_select_adj_719), 
            .debug_c_c(debug_c_c), .n30358(n30358), .\register_addr[0] (register_addr[0]), 
            .n30340(n30340), .n30406(n30406), .n30422(n30422), .n30445(n30445), 
            .rw(rw), .n30349(n30349), .n32380(n32380), .n9122(n9122), 
            .\quadA_delayed[1] (quadA_delayed_adj_1102[1]), .qreset(qreset), 
            .n6(n6_adj_603), .\quadB_delayed[1] (quadB_delayed_adj_1103[1]), 
            .n14013(n14013), .debug_c_0(debug_c_0), .encoder_li_c(encoder_li_c), 
            .encoder_lb_c(encoder_lb_c), .encoder_la_c(encoder_la_c), .\read_size[2] (read_size_adj_994[2]), 
            .n14291(n14291), .n30366(n30366), .read_value({read_value_adj_993}), 
            .\read_size[0] (read_size_adj_994[0]), .n302(n302), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(649[20] 659[47])
    LUT4 Select_4225_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[2]), 
         .D(rw), .Z(n8_adj_758)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4225_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4224_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[3]), 
         .D(rw), .Z(n8)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4224_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4150_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[31]), 
         .D(rw), .Z(n6_adj_755)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4150_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4153_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[30]), 
         .D(n32379), .Z(n6_adj_757)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4153_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i14295_3_lut (.A(Stepper_Z_En_c), .B(div_factor_reg_adj_909[6]), 
         .C(register_addr[1]), .Z(n20671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i14295_3_lut.init = 16'hcaca;
    \ClockDividerP_SP(factor=120000)  clk_100Hz_divider (.GND_net(GND_net), 
            .debug_c_0(debug_c_0), .debug_c_c(debug_c_c), .n32385(n32385), 
            .n32380(n32380)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(621[29] 623[61])
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .debug_c_c(debug_c_c), 
            .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_Z_nFault_c(Stepper_Z_nFault_c), 
            .n32382(n32382), .\read_size[0] (read_size_adj_912[0]), .n13918(n13918), 
            .n28323(n28323), .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n579(n571_adj_930[0]), 
            .prev_step_clk(prev_step_clk_adj_606), .step_clk(step_clk_adj_605), 
            .n13594(n13594), .prev_select(prev_select_adj_641), .n30391(n30391), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .n32(n32_adj_528), .n30422(n30422), 
            .\register_addr[2] (register_addr[2]), .n26507(n26507), .\register_addr[3] (register_addr[3]), 
            .n32380(n32380), .n26486(n26486), .read_value({read_value_adj_911}), 
            .\steps_reg[5] (steps_reg_adj_910[5]), .\steps_reg[6] (steps_reg_adj_910[6]), 
            .\steps_reg[9] (steps_reg_adj_910[9]), .\steps_reg[3] (steps_reg_adj_910[3]), 
            .databus({databus}), .n3892(n3892), .n13269(n13269), .\register_addr[4] (register_addr[4]), 
            .n30344(n30344), .\register_addr[5] (register_addr[5]), .limit_c_2(limit_c_2), 
            .n30421(n30421), .int_step(int_step), .n22(n22_adj_523), .n30310(n30310), 
            .n30317(n30317), .n32385(n32385), .n32381(n32381), .n32386(n32386), 
            .\div_factor_reg[9] (div_factor_reg_adj_909[9]), .\div_factor_reg[6] (div_factor_reg_adj_909[6]), 
            .\div_factor_reg[5] (div_factor_reg_adj_909[5]), .\div_factor_reg[3] (div_factor_reg_adj_909[3]), 
            .\control_reg[7] (control_reg_adj_908[7]), .Stepper_Z_En_c(Stepper_Z_En_c), 
            .Stepper_Z_Dir_c(Stepper_Z_Dir_c), .\control_reg[3] (control_reg_adj_908[3]), 
            .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), .\read_size[2] (read_size_adj_912[2]), 
            .n30342(n30342), .n20670(n20670), .n20681(n20681), .n6917(n6891[6]), 
            .n28148(n28148), .n8272(n8271[7])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(588[25] 601[45])
    LUT4 i14303_3_lut (.A(Stepper_Z_Dir_c), .B(div_factor_reg_adj_909[5]), 
         .C(register_addr[1]), .Z(n20679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i14303_3_lut.init = 16'hcaca;
    SabertoothSerialPeripheral motor_serial (.debug_c_c(debug_c_c), .n9122(n9122), 
            .n282(n281[15]), .n32384(n32384), .\databus[6] (databus[6]), 
            .\databus[5] (databus[5]), .\databus[4] (databus[4]), .\databus[3] (databus[3]), 
            .\databus[2] (databus[2]), .\databus[1] (databus[1]), .\databus[0] (databus[0]), 
            .n32385(n32385), .\read_size[0] (read_size_adj_852[0]), .n21563(n21563), 
            .n32381(n32381), .\select[2] (select[2]), .\register_addr[0] (register_addr[0]), 
            .n30422(n30422), .\register_addr[1] (register_addr[1]), .\register_addr[3] (register_addr[3]), 
            .\register_addr[2] (register_addr[2]), .n30445(n30445), .n32380(n32380), 
            .rw(rw), .n5(n5_adj_763), .n5_adj_221(n5), .n5_adj_222(n5_adj_766), 
            .n5_adj_223(n5_adj_759), .n5_adj_224(n5_adj_771), .n5_adj_225(n5_adj_769), 
            .n5_adj_226(n5_adj_773), .n5_adj_227(n5_adj_776), .n30488(n30488), 
            .n13269(n13269), .n30350(n30350), .n30314(n30314), .n30324(n30324), 
            .n13534(n13534), .n30349(n30349), .n30491(n30491), .n30489(n30489), 
            .n30379(n30379), .n28137(n28137), .n30478(n30478), .n8(n8_adj_681), 
            .\state[0] (state_adj_1038[0]), .GND_net(GND_net), .n12(n32520[0]), 
            .n30305(n30305), .n31(n31), .n27462(n27462), .n22(n22_adj_817), 
            .n19(n19_adj_827), .n32382(n32382), .\reset_count[14] (reset_count[14]), 
            .\reset_count[12] (reset_count[12]), .n28605(n28605), .motor_pwm_l_c(motor_pwm_l_c), 
            .n30342(n30342), .select_clk(select_clk), .n107(n107), .n8129(n8129)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(508[29] 516[56])
    LUT4 Select_4156_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[29]), 
         .D(n32379), .Z(n6_adj_756)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4156_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4159_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[28]), 
         .D(n32379), .Z(n6_adj_563)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4159_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4162_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[27]), 
         .D(n32379), .Z(n6_adj_810)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4162_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i14292_3_lut (.A(control_reg_adj_908[3]), .B(div_factor_reg_adj_909[3]), 
         .C(register_addr[1]), .Z(n20668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i14292_3_lut.init = 16'hcaca;
    LUT4 Select_4165_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[26]), 
         .D(n32379), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4165_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4168_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[25]), 
         .D(rw), .Z(n6_adj_812)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4168_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    \ProtocolInterface(baud_div=12)  protocol_interface (.register_addr({Open_0, 
            Open_1, register_addr[5:2], Open_2, register_addr[0]}), 
            .debug_c_c(debug_c_c), .databus({databus}), .debug_c_5(debug_c_5), 
            .\select[4] (select[4]), .n30491(n30491), .n30489(n30489), 
            .n30479(n30479), .n30391(n30391), .n30488(n30488), .n30396(n30396), 
            .n30398(n30398), .sendcount({Open_3, Open_4, Open_5, Open_6, 
            sendcount[0]}), .n13574(n13574), .databus_out({databus_out}), 
            .n32377(n32377), .n32379(n32379), .prev_select(prev_select_adj_678), 
            .\read_value[1] (read_value_adj_952[1]), .rw(rw), .n1(n1_adj_761), 
            .n32380(n32380), .n2673(n2673), .\select[7] (select[7]), .\sendcount[3] (sendcount[3]), 
            .\select[3] (select[3]), .\select[2] (select[2]), .\select[1] (select[1]), 
            .debug_c_7(debug_c_7), .n30383(n30383), .n3806(n3806), .n5632(n5632), 
            .n26671(n26671), .n32376(n32376), .n30321(n30321), .\register[1][0] (\register[1]_adj_1000 [0]), 
            .n97(n99_adj_1268[0]), .\register[1][24] (\register[1]_adj_1000 [24]), 
            .n49(n99_adj_1268[24]), .n1307(n1295[20]), .n28421(n28421), 
            .n1313(n1295[14]), .n1310(n1295[17]), .\register[1][25] (\register[1]_adj_1000 [25]), 
            .n47(n99_adj_1268[25]), .\register[1][29] (\register[1]_adj_1000 [29]), 
            .n39(n99_adj_1268[29]), .n30316(n30316), .n3666(n3666), .debug_c_2(debug_c_2), 
            .debug_c_3(debug_c_3), .\register[1][30] (\register[1]_adj_1000 [30]), 
            .n37(n99_adj_1268[30]), .debug_c_4(debug_c_4), .n30324(n30324), 
            .n21310(n21310), .n3989(n3989), .n30344(n30344), .n3892(n3892), 
            .n30422(n30422), .\register_addr[1] (register_addr[1]), .n30411(n30411), 
            .n30394(n30394), .n30413(n30413), .n30385(n30385), .n17(n17_adj_525), 
            .n4(n4_adj_820), .\reg_size[2] (reg_size[2]), .n30454(n30454), 
            .\steps_reg[7] (steps_reg_adj_951[7]), .n19(n19_adj_679), .\control_reg[7] (control_reg[7]), 
            .n1_adj_216(n1), .\steps_reg[4] (steps_reg_adj_869[4]), .n17_adj_217(n17), 
            .n4_adj_218(n4_adj_821), .\steps_reg[6] (steps_reg_adj_910[6]), 
            .n13(n13), .n30373(n30373), .n30417(n30417), .n28218(n28218), 
            .n30317(n30317), .\steps_reg[5] (steps_reg_adj_910[5]), .n14(n14), 
            .\steps_reg[3] (steps_reg_adj_910[3]), .n12(n12), .\control_reg[7]_adj_219 (control_reg_adj_867[7]), 
            .n8263(n8262[7]), .\control_reg[7]_adj_220 (control_reg_adj_908[7]), 
            .n8272(n8271[7]), .\reset_count[14] (reset_count[14]), .\reset_count[13] (reset_count[13]), 
            .\reset_count[12] (reset_count[12]), .n26787(n26787), .n10643(n10643), 
            .GND_net(GND_net), .uart_rx_c(uart_rx_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[26] 485[57])
    LUT4 Select_4171_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[24]), 
         .D(rw), .Z(n6_adj_808)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4171_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4174_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[23]), 
         .D(rw), .Z(n6_adj_818)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4174_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4177_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[22]), 
         .D(n32379), .Z(n6_adj_806)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4177_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4180_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[21]), 
         .D(rw), .Z(n6_adj_797)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4180_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4183_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[20]), 
         .D(rw), .Z(n6_adj_795)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4183_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4186_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[19]), 
         .D(rw), .Z(n6_adj_799)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4186_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 Select_4189_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[18]), 
         .D(rw), .Z(n6_adj_796)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4189_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 m1_lut (.Z(n32376)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.debug_c_c(debug_c_c), .n8894(n8894), 
            .n32384(n32384), .databus({databus}), .n608(n580[4]), .n610(n580_adj_890[2]), 
            .\control_reg[7] (control_reg_adj_867[7]), .Stepper_Y_En_c(Stepper_Y_En_c), 
            .Stepper_Y_Dir_c(Stepper_Y_Dir_c), .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), 
            .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), .\read_size[2] (read_size_adj_871[2]), 
            .n14121(n14121), .\steps_reg[24] (steps_reg_adj_869[24]), .n32385(n32385), 
            .n32381(n32381), .n32382(n32382), .\steps_reg[20] (steps_reg_adj_869[20]), 
            .n3666(n3666), .n32383(n32383), .\steps_reg[4] (steps_reg_adj_869[4]), 
            .\steps_reg[1] (steps_reg_adj_869[1]), .\register_addr[1] (register_addr[1]), 
            .fault_latched(fault_latched), .VCC_net(VCC_net), .GND_net(GND_net), 
            .Stepper_Y_nFault_c(Stepper_Y_nFault_c), .\read_size[0] (read_size_adj_871[0]), 
            .n32(n32), .\register_addr[2] (register_addr[2]), .\register_addr[3] (register_addr[3]), 
            .\register_addr[4] (register_addr[4]), .n28196(n28196), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), 
            .n579(n571_adj_930[0]), .prev_step_clk(prev_step_clk_adj_566), 
            .step_clk(step_clk_adj_565), .prev_select(prev_select_adj_601), 
            .n30374(n30374), .read_value({read_value_adj_870}), .n9128(n9128), 
            .n26485(n26485), .\register_addr[0] (register_addr[0]), .n30370(n30370), 
            .n30380(n30380), .n30421(n30421), .\register_addr[5] (register_addr[5]), 
            .limit_c_1(limit_c_1), .Stepper_Y_Step_c(Stepper_Y_Step_c), 
            .n30489(n30489), .n30491(n30491), .\select[4] (select[4]), 
            .n30427(n30427), .n30406(n30406), .n30417(n30417), .n28184(n28184), 
            .n32380(n32380), .n30316(n30316), .n13269(n13269), .n30331(n30331), 
            .rw(rw), .n22(n22), .n30311(n30311), .n21533(n21533), .n28324(n28324), 
            .n30479(n30479), .n28323(n28323), .n12(n12_adj_642), .n28172(n28172), 
            .n19585(n19585), .n30342(n30342), .\div_factor_reg[24] (div_factor_reg_adj_868[24]), 
            .n28672(n28672), .\div_factor_reg[1] (div_factor_reg_adj_868[1]), 
            .n49(n99_adj_1273[24]), .\div_factor_reg[20] (div_factor_reg_adj_868[20]), 
            .n17(n17), .n8263(n8262[7])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(573[25] 586[45])
    PFUMX i14305 (.BLUT(n20679), .ALUT(n14), .C0(register_addr[0]), .Z(n20681));
    LUT4 i21698_2_lut (.A(n28748), .B(n32380), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21698_2_lut.init = 16'heeee;
    ClockDivider_U10 pwm_clk_div (.debug_c_c(debug_c_c), .n241(n241), .n32380(n32380), 
            .n7504(n7504), .n30303(n30303), .n28775(n28775), .n26601(n26601), 
            .n28723(n28723), .n26592(n26592), .GND_net(GND_net), .n28725(n28725), 
            .n26596(n26596), .n28910(n28910), .n13624(n13624), .n28859(n28859), 
            .n14284(n14284), .n28857(n28857), .n14306(n14306), .n28855(n28855), 
            .n14307(n14307), .n28853(n28853), .n14308(n14308), .n28851(n28851), 
            .n14309(n14309), .n28765(n28765), .n26618(n26618), .n28770(n28770), 
            .n26607(n26607), .n28773(n28773), .n26604(n26604)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(518[15] 521[41])
    LUT4 Select_4192_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n30385), .C(read_value_adj_1002[17]), 
         .D(rw), .Z(n6_adj_805)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(631[4] 647[11])
    defparam Select_4192_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21696_4_lut (.A(n13_adj_814), .B(n30444), .C(n11_adj_815), .D(n20944), 
         .Z(n28748)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21696_4_lut.init = 16'h0001;
    LUT4 i5_4_lut (.A(reset_count[5]), .B(reset_count[12]), .C(reset_count[0]), 
         .D(reset_count[1]), .Z(n13_adj_814)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(reset_count[3]), .B(reset_count[2]), .Z(n11_adj_815)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam i3_2_lut.init = 16'heeee;
    RCPeripheral rc_receiver (.read_value({read_value}), .\read_value[7]_adj_7 (read_value_adj_870[7]), 
            .n46(n46), .n3(n3_adj_783), .databus({databus}), .\read_value[13]_adj_8 (read_value_adj_952[13]), 
            .read_value_adj_215({read_value_adj_993}), .n47(n47), .\read_value[7]_adj_41 (read_value_adj_858[7]), 
            .n30372(n30372), .\read_value[13]_adj_42 (read_value_adj_858[13]), 
            .n6(n6_adj_785), .databus_out({databus_out}), .n32379(n32379), 
            .n8(n8_adj_767), .\register_addr[0] (register_addr[0]), .\register_addr[1] (register_addr[1]), 
            .n3_adj_43(n3_adj_680), .\select[7] (select[7]), .n30395(n30395), 
            .n176(n176), .n2(n2_adj_770), .\read_value[5]_adj_44 (read_value_adj_870[5]), 
            .n3_adj_45(n3_adj_782), .\read_value[11]_adj_46 (read_value_adj_952[11]), 
            .\read_value[11]_adj_47 (read_value_adj_858[11]), .n6_adj_48(n6_adj_784), 
            .\read_value[11]_adj_49 (read_value_adj_911[11]), .n30367(n30367), 
            .\read_value[26]_adj_50 (read_value_adj_952[26]), .read_size({read_size}), 
            .\select[1] (select[1]), .n30454(n30454), .\reg_size[2] (reg_size[2]), 
            .\sendcount[3] (sendcount[3]), .n4(n4_adj_820), .n3_adj_51(n3_adj_823), 
            .\read_value[13]_adj_52 (read_value_adj_911[13]), .\read_value[31]_adj_53 (read_value_adj_952[31]), 
            .\register_addr[4] (register_addr[4]), .n30427(n30427), .\register_addr[5] (register_addr[5]), 
            .n30371(n30371), .\read_value[31]_adj_54 (read_value_adj_858[31]), 
            .n6_adj_55(n6_adj_755), .rw(rw), .\read_value[31]_adj_56 (read_value_adj_911[31]), 
            .\read_value[6]_adj_57 (read_value_adj_952[6]), .n5(n5_adj_773), 
            .prev_select(prev_select_adj_678), .n32377(n32377), .n30338(n30338), 
            .n30374(n30374), .prev_select_adj_58(prev_select_adj_601), .n30331(n30331), 
            .n3_adj_59(n3_adj_778), .\read_value[10]_adj_60 (read_value_adj_952[10]), 
            .\read_value[10]_adj_61 (read_value_adj_858[10]), .n6_adj_62(n6_adj_780), 
            .n3_adj_63(n3_adj_822), .\read_value[30]_adj_64 (read_value_adj_952[30]), 
            .\read_value[30]_adj_65 (read_value_adj_858[30]), .n6_adj_66(n6_adj_757), 
            .\read_value[30]_adj_67 (read_value_adj_911[30]), .n3_adj_68(n3_adj_524), 
            .\read_value[29]_adj_69 (read_value_adj_952[29]), .\read_value[29]_adj_70 (read_value_adj_858[29]), 
            .n6_adj_71(n6_adj_756), .\read_value[10]_adj_72 (read_value_adj_911[10]), 
            .\read_value[29]_adj_73 (read_value_adj_911[29]), .n3_adj_74(n3_adj_602), 
            .\read_value[28]_adj_75 (read_value_adj_952[28]), .\read_value[28]_adj_76 (read_value_adj_858[28]), 
            .n6_adj_77(n6_adj_563), .\read_value[28]_adj_78 (read_value_adj_911[28]), 
            .n8_adj_79(n8_adj_774), .\read_value[6]_adj_80 (read_value_adj_870[6]), 
            .n3_adj_81(n3_adj_809), .\read_value[6]_adj_82 (read_value_adj_858[6]), 
            .\read_value[27]_adj_83 (read_value_adj_952[27]), .n3_adj_84(n3_adj_788), 
            .\read_value[27]_adj_85 (read_value_adj_858[27]), .n6_adj_86(n6_adj_810), 
            .\read_value[27]_adj_87 (read_value_adj_911[27]), .\read_value[5]_adj_88 (read_value_adj_952[5]), 
            .n5_adj_89(n5_adj_769), .n2_adj_90(n2_adj_768), .\read_value[5]_adj_91 (read_value_adj_858[5]), 
            .\read_value[26]_adj_92 (read_value_adj_858[26]), .n6_adj_93(n6), 
            .\read_value[9]_adj_94 (read_value_adj_952[9]), .\read_value[26]_adj_95 (read_value_adj_911[26]), 
            .n3_adj_96(n3_adj_811), .\read_value[25]_adj_97 (read_value_adj_952[25]), 
            .\read_value[9]_adj_98 (read_value_adj_858[9]), .n6_adj_99(n6_adj_789), 
            .\register_addr[2] (register_addr[2]), .\read_value[9]_adj_100 (read_value_adj_911[9]), 
            .n2_adj_101(n2_adj_775), .\read_value[7]_adj_102 (read_value_adj_952[7]), 
            .n5_adj_103(n5_adj_776), .n8_adj_104(n8_adj_777), .\read_value[25]_adj_105 (read_value_adj_858[25]), 
            .n6_adj_106(n6_adj_812), .\read_value[25]_adj_107 (read_value_adj_911[25]), 
            .n3_adj_108(n3_adj_807), .n2_adj_109(n2_adj_826), .\read_value[24]_adj_110 (read_value_adj_952[24]), 
            .\read_value[24]_adj_111 (read_value_adj_858[24]), .n6_adj_112(n6_adj_808), 
            .n2_adj_113(n2_adj_764), .\read_value[24]_adj_114 (read_value_adj_911[24]), 
            .\read_value[0]_adj_115 (read_value_adj_952[0]), .n5_adj_116(n5_adj_763), 
            .n3_adj_117(n3_adj_813), .\read_value[4]_adj_118 (read_value_adj_952[4]), 
            .n5_adj_119(n5_adj_771), .n8_adj_120(n8_adj_772), .\read_value[23]_adj_121 (read_value_adj_952[23]), 
            .\read_value[4]_adj_122 (read_value_adj_870[4]), .\read_value[23]_adj_123 (read_value_adj_858[23]), 
            .n6_adj_124(n6_adj_818), .\read_value[23]_adj_125 (read_value_adj_911[23]), 
            .n2_adj_126(n2_adj_760), .n3_adj_127(n3_adj_800), .\read_value[4]_adj_128 (read_value_adj_858[4]), 
            .\read_value[22]_adj_129 (read_value_adj_952[22]), .\read_value[22]_adj_130 (read_value_adj_858[22]), 
            .n6_adj_131(n6_adj_806), .\read_value[22]_adj_132 (read_value_adj_911[22]), 
            .n3_adj_133(n3), .\read_value[21]_adj_134 (read_value_adj_952[21]), 
            .\read_value[21]_adj_135 (read_value_adj_858[21]), .n6_adj_136(n6_adj_797), 
            .n8_adj_137(n8_adj_762), .\read_value[21]_adj_138 (read_value_adj_911[21]), 
            .n3_adj_139(n3_adj_801), .\read_value[20]_adj_140 (read_value_adj_952[20]), 
            .\read_value[20]_adj_141 (read_value_adj_858[20]), .n6_adj_142(n6_adj_795), 
            .\read_value[20]_adj_143 (read_value_adj_911[20]), .n3_adj_144(n3_adj_798), 
            .\read_value[19]_adj_145 (read_value_adj_952[19]), .\read_value[19]_adj_146 (read_value_adj_858[19]), 
            .n6_adj_147(n6_adj_799), .\read_value[19]_adj_148 (read_value_adj_911[19]), 
            .n3_adj_149(n3_adj_794), .\read_value[18]_adj_150 (read_value_adj_952[18]), 
            .\read_value[18]_adj_151 (read_value_adj_858[18]), .n6_adj_152(n6_adj_796), 
            .\read_value[18]_adj_153 (read_value_adj_911[18]), .n3_adj_154(n3_adj_804), 
            .\read_value[17]_adj_155 (read_value_adj_952[17]), .\read_value[17]_adj_156 (read_value_adj_858[17]), 
            .n6_adj_157(n6_adj_805), .\read_value[17]_adj_158 (read_value_adj_911[17]), 
            .n3_adj_159(n3_adj_802), .\read_value[16]_adj_160 (read_value_adj_952[16]), 
            .\read_value[16]_adj_161 (read_value_adj_858[16]), .n6_adj_162(n6_adj_803), 
            .\read_value[16]_adj_163 (read_value_adj_911[16]), .n3_adj_164(n3_adj_792), 
            .\read_value[15]_adj_165 (read_value_adj_952[15]), .\read_value[15]_adj_166 (read_value_adj_858[15]), 
            .n6_adj_167(n6_adj_793), .\read_value[15]_adj_168 (read_value_adj_911[15]), 
            .n3_adj_169(n3_adj_790), .\read_value[14]_adj_170 (read_value_adj_952[14]), 
            .\read_value[14]_adj_171 (read_value_adj_858[14]), .n6_adj_172(n6_adj_791), 
            .\read_value[14]_adj_173 (read_value_adj_911[14]), .n2_adj_174(n2), 
            .\read_value[2]_adj_175 (read_value_adj_952[2]), .n5_adj_176(n5_adj_759), 
            .n3_adj_177(n3_adj_779), .\read_value[12]_adj_178 (read_value_adj_952[12]), 
            .\read_value[12]_adj_179 (read_value_adj_858[12]), .n6_adj_180(n6_adj_781), 
            .\read_value[12]_adj_181 (read_value_adj_911[12]), .n8_adj_182(n8_adj_758), 
            .n3_adj_183(n3_adj_786), .\read_value[8]_adj_184 (read_value_adj_952[8]), 
            .\read_value[8]_adj_185 (read_value_adj_858[8]), .n6_adj_186(n6_adj_787), 
            .\read_value[8]_adj_187 (read_value_adj_911[8]), .\read_size[0]_adj_188 (read_size_adj_1003[0]), 
            .n30361(n30361), .n11(n11), .n30396(n30396), .\read_size[0]_adj_189 (read_size_adj_859[0]), 
            .n16(n16_adj_682), .\read_size[0]_adj_190 (read_size_adj_953[0]), 
            .\read_size[0]_adj_191 (read_size_adj_994[0]), .n30358(n30358), 
            .n12(n12_adj_683), .\read_size[0]_adj_192 (read_size_adj_871[0]), 
            .\read_size[0]_adj_193 (read_size_adj_912[0]), .\read_size[0]_adj_194 (read_size_adj_852[0]), 
            .n30391(n30391), .\select[2] (select[2]), .\read_size[2]_adj_195 (read_size_adj_1003[2]), 
            .\read_value[0]_adj_196 (read_value_adj_870[0]), .\read_size[2]_adj_197 (read_size_adj_994[2]), 
            .\read_value[1]_adj_198 (read_value_adj_870[1]), .\read_value[2]_adj_199 (read_value_adj_870[2]), 
            .n4_adj_200(n4), .\read_value[2]_adj_201 (read_value_adj_858[2]), 
            .\read_value[0]_adj_202 (read_value_adj_858[0]), .\read_value[1]_adj_203 (read_value_adj_1002[1]), 
            .n30339(n30339), .n2_adj_204(n2_adj_765), .\read_size[2]_adj_205 (read_size_adj_859[2]), 
            .\read_size[2]_adj_206 (read_size_adj_871[2]), .\read_size[2]_adj_207 (read_size_adj_912[2]), 
            .\read_size[2]_adj_208 (read_size_adj_953[2]), .\read_value[3]_adj_209 (read_value_adj_952[3]), 
            .n5_adj_210(n5_adj_766), .n8_adj_211(n8), .\read_value[3]_adj_212 (read_value_adj_870[3]), 
            .\read_value[3]_adj_213 (read_value_adj_858[3]), .n1(n1_adj_761), 
            .n5_adj_214(n5), .GND_net(GND_net), .n28765(n28765), .debug_c_c(debug_c_c), 
            .n30303(n30303), .rc_ch8_c(rc_ch8_c), .n26618(n26618), .n28910(n28910), 
            .n13624(n13624), .rc_ch7_c(rc_ch7_c), .n26601(n26601), .n28859(n28859), 
            .n28775(n28775), .n14284(n14284), .rc_ch4_c(rc_ch4_c), .n28857(n28857), 
            .n14306(n14306), .n28723(n28723), .n26592(n26592), .n28855(n28855), 
            .rc_ch3_c(rc_ch3_c), .n26607(n26607), .n14307(n14307), .n28770(n28770), 
            .n28853(n28853), .n26604(n26604), .n14308(n14308), .rc_ch2_c(rc_ch2_c), 
            .n28773(n28773), .n32380(n32380), .n28851(n28851), .n14309(n14309), 
            .rc_ch1_c(rc_ch1_c), .n28725(n28725), .n26596(n26596)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(673[15] 685[41])
    EncoderPeripheral right_encoder (.read_value({read_value_adj_1002}), .debug_c_c(debug_c_c), 
            .n13589(n13589), .n30321(n30321), .\read_size[2] (read_size_adj_1003[2]), 
            .n30380(n30380), .\register_addr[0] (register_addr[0]), .\read_size[0] (read_size_adj_1003[0]), 
            .n30370(n30370), .prev_select(prev_select_adj_754), .n30361(n30361), 
            .encoder_ra_c(encoder_ra_c), .encoder_rb_c(encoder_rb_c), .encoder_ri_c(encoder_ri_c), 
            .\register_addr[1] (register_addr[1]), .n30489(n30489), .n30491(n30491), 
            .n13269(n13269), .n30422(n30422), .n30366(n30366), .n302(n302), 
            .n97(n99_adj_1268[0]), .n49(n99_adj_1268[24]), .n47(n99_adj_1268[25]), 
            .n39(n99_adj_1268[29]), .n37(n99_adj_1268[30]), .n14013(n14013), 
            .qreset(qreset), .\quadA_delayed[1] (quadA_delayed_adj_1102[1]), 
            .GND_net(GND_net), .n6(n6_adj_603), .\register[1][0] (\register[1]_adj_1000 [0]), 
            .VCC_net(VCC_net), .\register[1][24] (\register[1]_adj_1000 [24]), 
            .\register[1][25] (\register[1]_adj_1000 [25]), .\register[1][29] (\register[1]_adj_1000 [29]), 
            .\register[1][30] (\register[1]_adj_1000 [30]), .\quadB_delayed[1] (quadB_delayed_adj_1103[1])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(660[20] 670[47])
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.debug_c_c(debug_c_c), .n8890(n8890), 
            .n32383(n32383), .databus({databus}), .n608(n580[4]), .n610(n580_adj_890[2]), 
            .\control_reg[7] (control_reg[7]), .n30314(n30314), .Stepper_X_En_c(Stepper_X_En_c), 
            .Stepper_X_Dir_c(Stepper_X_Dir_c), .n13534(n13534), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\read_size[2] (read_size_adj_859[2]), 
            .n2644(n2644), .n28137(n28137), .n32384(n32384), .n32381(n32381), 
            .n32382(n32382), .\read_size[0] (read_size_adj_859[0]), .n21563(n21563), 
            .Stepper_X_M0_c_0(Stepper_X_M0_c_0), .n579(n571_adj_930[0]), 
            .prev_step_clk(prev_step_clk), .step_clk(step_clk), .prev_select(prev_select), 
            .n30396(n30396), .read_value({read_value_adj_858}), .n9125(n9125), 
            .\register_addr[1] (register_addr[1]), .n11(n11_adj_816), .\register_addr[0] (register_addr[0]), 
            .n30330(n30330), .n3989(n3989), .n30422(n30422), .n30307(n30307), 
            .n30489(n30489), .n28421(n28421), .n9118(n9118), .limit_c_0(limit_c_0), 
            .Stepper_X_Step_c(Stepper_X_Step_c), .n34(n34), .n26484(n26484), 
            .n24(n24), .n30313(n30313), .n1(n1), .GND_net(GND_net), 
            .VCC_net(VCC_net), .Stepper_X_nFault_c(Stepper_X_nFault_c), 
            .n32380(n32380), .n32385(n32385)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(558[25] 571[45])
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.read_value({read_value_adj_952}), 
            .debug_c_c(debug_c_c), .n2673(n2673), .n9136(n9136), .n32382(n32382), 
            .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_953[0]), .n28324(n28324), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .databus({databus}), .prev_select(prev_select_adj_678), .n30371(n30371), 
            .n32383(n32383), .n32381(n32381), .\control_reg[7] (control_reg_adj_949[7]), 
            .Stepper_A_En_c(Stepper_A_En_c), .Stepper_A_Dir_c(Stepper_A_Dir_c), 
            .Stepper_A_M2_c_2(Stepper_A_M2_c_2), .Stepper_A_M1_c_1(Stepper_A_M1_c_1), 
            .\register_addr[0] (register_addr[0]), .n3806(n3806), .\register_addr[1] (register_addr[1]), 
            .stepping(stepping), .n26585(n26585), .\steps_reg[7] (steps_reg_adj_951[7]), 
            .\register_addr[5] (register_addr[5]), .\register_addr[4] (register_addr[4]), 
            .n21533(n21533), .limit_c_3(limit_c_3), .Stepper_A_Step_c(Stepper_A_Step_c), 
            .n30491(n30491), .n28218(n28218), .rw(rw), .n30338(n30338), 
            .n13269(n13269), .n28184(n28184), .n30411(n30411), .n32380(n32380), 
            .\read_size[2] (read_size_adj_953[2]), .n28172(n28172), .n32(n32_adj_528), 
            .prev_step_clk(prev_step_clk_adj_606), .step_clk(step_clk_adj_605), 
            .n30310(n30310), .n32385(n32385), .n32386(n32386), .n22(n22_adj_523), 
            .n32_adj_1(n32), .prev_step_clk_adj_2(prev_step_clk_adj_566), 
            .step_clk_adj_3(step_clk_adj_565), .n30311(n30311), .n22_adj_4(n22), 
            .prev_step_clk_adj_5(prev_step_clk), .n34(n34), .step_clk_adj_6(step_clk), 
            .n30313(n30313), .n24(n24), .n19(n19_adj_679)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(603[25] 616[45])
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (debug_c_c, n32384, \databus[1] , \select[1] , 
            rw, n46, n32381, read_size, n30307, n302, n26507, 
            n30330, n32380, n32385, \register_addr[4] , \register_addr[3] , 
            n21310, xbee_pause_c, \register_addr[0] , n9118, n30478, 
            n11, \register_addr[1] , n30366, n30413, \register_addr[2] , 
            n6, n30491, n28421, n30395, n176, n8, \control_reg[7] , 
            n26486, n32, \control_reg[7]_adj_228 , n26485, n32_adj_229, 
            \control_reg[7]_adj_230 , n26585, stepping, \control_reg[7]_adj_231 , 
            n26484, n34, \state[0] , n22, n27462, signal_light_c, 
            n31, n19, n28218, n30344, n30417, n13594, n32377, 
            \select[3] , n30358, \register_addr[5] , n30361, read_value, 
            GND_net, n30394, n30324, n30489, n8890) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n32384;
    input \databus[1] ;
    input \select[1] ;
    input rw;
    output n46;
    input n32381;
    output [2:0]read_size;
    output n30307;
    input n302;
    input n26507;
    input n30330;
    input n32380;
    input n32385;
    input \register_addr[4] ;
    input \register_addr[3] ;
    output n21310;
    input xbee_pause_c;
    input \register_addr[0] ;
    input n9118;
    output n30478;
    output n11;
    input \register_addr[1] ;
    input n30366;
    input n30413;
    input \register_addr[2] ;
    input n6;
    input n30491;
    input n28421;
    output n30395;
    output n176;
    input n8;
    input \control_reg[7] ;
    input n26486;
    output n32;
    input \control_reg[7]_adj_228 ;
    input n26485;
    output n32_adj_229;
    input \control_reg[7]_adj_230 ;
    input n26585;
    output stepping;
    input \control_reg[7]_adj_231 ;
    input n26484;
    output n34;
    input \state[0] ;
    input n22;
    output n27462;
    output signal_light_c;
    input n31;
    output n19;
    input n28218;
    input n30344;
    input n30417;
    output n13594;
    input n32377;
    input \select[3] ;
    output n30358;
    input \register_addr[5] ;
    output n30361;
    output [31:0]read_value;
    input GND_net;
    input n30394;
    input n30324;
    input n30489;
    output n8890;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire force_pause, n26278;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n13814;
    wire [31:0]n100;
    
    wire prev_clk_1Hz, clk_1Hz;
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n178, prev_select;
    wire [31:0]n5772;
    
    wire n30433, n28052;
    wire [31:0]n99;
    
    wire n30475, n16115, n16116, n29649, n21215, n26670, n25814, 
        n25813, n25812, n25811, n25810, n25809, n25808, n28599, 
        n25807, n25806, n25805, n25804, n25803, n25802, n25801, 
        n25800, n25799, n29650, n29613, n29612;
    
    FD1P3IX force_pause_151 (.D(\databus[1] ), .SP(n26278), .CD(n32384), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam force_pause_151.GSR = "ENABLED";
    LUT4 i14_2_lut (.A(\select[1] ), .B(rw), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam i14_2_lut.init = 16'h8888;
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n13814), .CD(n32381), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n302), .SP(n30307), .CK(debug_c_c), .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_149 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_clk_1Hz_149.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_150 (.D(n178), .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam xbee_pause_latched_150.GSR = "ENABLED";
    FD1S3AX prev_select_148 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_select_148.GSR = "ENABLED";
    LUT4 i14930_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [22]), 
         .Z(n5772[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14930_2_lut_3_lut.init = 16'h2020;
    LUT4 i134_2_lut_rep_424 (.A(prev_clk_1Hz), .B(clk_1Hz), .Z(n30433)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i134_2_lut_rep_424.init = 16'h4444;
    LUT4 i14927_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [23]), 
         .Z(n5772[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14927_2_lut_3_lut.init = 16'h2020;
    LUT4 i14926_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [24]), 
         .Z(n5772[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14926_2_lut_3_lut.init = 16'h2020;
    LUT4 i14925_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [25]), 
         .Z(n5772[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14925_2_lut_3_lut.init = 16'h2020;
    LUT4 i2695_2_lut_3_lut (.A(prev_clk_1Hz), .B(clk_1Hz), .C(n32380), 
         .Z(n13814)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i2695_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i14920_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [26]), 
         .Z(n5772[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14920_2_lut_3_lut.init = 16'h2020;
    LUT4 i14919_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [27]), 
         .Z(n5772[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14919_2_lut_3_lut.init = 16'h2020;
    LUT4 i14918_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [28]), 
         .Z(n5772[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14918_2_lut_3_lut.init = 16'h2020;
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n30433), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n30433), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n13814), .CD(n32384), 
            .CK(debug_c_c), .Q(\register[2] [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n13814), .CD(n32384), 
            .CK(debug_c_c), .Q(\register[2] [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n13814), .CD(n32384), 
            .CK(debug_c_c), .Q(\register[2] [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n13814), .CD(n32384), 
            .CK(debug_c_c), .Q(\register[2] [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n13814), .CD(n32385), 
            .CK(debug_c_c), .Q(\register[2] [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    LUT4 i14897_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [29]), 
         .Z(n5772[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14897_2_lut_3_lut.init = 16'h2020;
    LUT4 i15124_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [30]), 
         .Z(n5772[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15124_2_lut_3_lut.init = 16'h2020;
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n13814), .CD(n32385), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    LUT4 i15125_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [31]), 
         .Z(n5772[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15125_2_lut_3_lut.init = 16'h2020;
    LUT4 i14935_2_lut (.A(\register_addr[4] ), .B(\register_addr[3] ), .Z(n21310)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14935_2_lut.init = 16'heeee;
    LUT4 i114_1_lut (.A(xbee_pause_c), .Z(n178)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(54[26:39])
    defparam i114_1_lut.init = 16'h5555;
    LUT4 i14835_4_lut (.A(\register_addr[0] ), .B(n9118), .C(n26507), 
         .D(n28052), .Z(n99[0])) /* synthesis lut_function=(!(A (B+(C))+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam i14835_4_lut.init = 16'h1303;
    LUT4 i1_4_lut (.A(n30478), .B(n11), .C(\register[2] [0]), .D(\register_addr[1] ), 
         .Z(n28052)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h3022;
    LUT4 i2_4_lut (.A(n32380), .B(rw), .C(n30475), .D(n30366), .Z(n26278)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam i2_4_lut.init = 16'h0032;
    LUT4 i3_3_lut_4_lut (.A(\register_addr[3] ), .B(n30413), .C(\register_addr[2] ), 
         .D(\register_addr[4] ), .Z(n11)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_rep_386 (.A(\register_addr[2] ), .B(n6), .C(n30491), 
         .D(n28421), .Z(n30395)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_rep_386.init = 16'hfefc;
    LUT4 i15295_1_lut_4_lut (.A(\register_addr[2] ), .B(n6), .C(n30491), 
         .D(n28421), .Z(n176)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+(C)))) */ ;
    defparam i15295_1_lut_4_lut.init = 16'h0103;
    LUT4 i117_2_lut_rep_466 (.A(prev_select), .B(\select[1] ), .Z(n30475)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i117_2_lut_rep_466.init = 16'h4444;
    LUT4 i9703_2_lut_3_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(n8), .D(n32380), .Z(n16115)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i9703_2_lut_3_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i9704_2_lut_3_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(n8), .D(n32380), .Z(n16116)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i9704_2_lut_3_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i947_2_lut_rep_298_2_lut_3_lut (.A(prev_select), .B(\select[1] ), 
         .C(n32380), .Z(n30307)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i947_2_lut_rep_298_2_lut_3_lut.init = 16'h0404;
    LUT4 i112_2_lut_rep_469 (.A(\register[0] [2]), .B(force_pause), .Z(n30478)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i112_2_lut_rep_469.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(\control_reg[7] ), 
         .D(n26486), .Z(n32)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_453 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_228 ), .D(n26485), .Z(n32_adj_229)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_453.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_454 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_230 ), .D(n26585), .Z(stepping)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_454.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_455 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_231 ), .D(n26484), .Z(n34)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_455.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_456 (.A(\register[0] [2]), .B(force_pause), 
         .C(\state[0] ), .D(n22), .Z(n27462)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_456.init = 16'h0100;
    LUT4 i14497_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(clk_1Hz), 
         .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i14497_2_lut_3_lut.init = 16'hfefe;
    LUT4 i21778_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(n31), 
         .D(\state[0] ), .Z(n19)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i21778_3_lut_4_lut.init = 16'h00ef;
    LUT4 i1_2_lut_4_lut (.A(n28218), .B(n30344), .C(n30417), .D(n32380), 
         .Z(n13594)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(64[8] 95[15])
    defparam i1_2_lut_4_lut.init = 16'hff80;
    LUT4 i14949_2_lut_rep_349_3_lut_4_lut (.A(n32377), .B(n30491), .C(\select[3] ), 
         .D(\register_addr[4] ), .Z(n30358)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i14949_2_lut_rep_349_3_lut_4_lut.init = 16'he0f0;
    LUT4 i14769_2_lut_rep_352_3_lut_4_lut (.A(\register_addr[5] ), .B(n30491), 
         .C(\select[3] ), .D(\register_addr[4] ), .Z(n30361)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i14769_2_lut_rep_352_3_lut_4_lut.init = 16'h1000;
    FD1P3AX read_value__i0 (.D(n99[0]), .SP(n30307), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 register_addr_0__bdd_4_lut (.A(\register_addr[0] ), .B(force_pause), 
         .C(\register_addr[1] ), .D(\register[2] [1]), .Z(n29649)) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam register_addr_0__bdd_4_lut.init = 16'h5e0e;
    LUT4 i14790_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [7]), 
         .Z(n5772[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14790_2_lut_3_lut.init = 16'h2020;
    LUT4 i21717_4_lut (.A(n30413), .B(n21310), .C(\register_addr[2] ), 
         .D(n21215), .Z(n26670)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i21717_4_lut.init = 16'h0111;
    LUT4 i14840_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n21215)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14840_2_lut.init = 16'heeee;
    CCU2D add_134_33 (.A0(\register[2] [31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25814), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_33.INIT0 = 16'h5aaa;
    defparam add_134_33.INIT1 = 16'h0000;
    defparam add_134_33.INJECT1_0 = "NO";
    defparam add_134_33.INJECT1_1 = "NO";
    CCU2D add_134_31 (.A0(\register[2] [29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25813), .COUT(n25814), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_31.INIT0 = 16'h5aaa;
    defparam add_134_31.INIT1 = 16'h5aaa;
    defparam add_134_31.INJECT1_0 = "NO";
    defparam add_134_31.INJECT1_1 = "NO";
    LUT4 i14548_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [15]), 
         .Z(n5772[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14548_2_lut_3_lut.init = 16'h2020;
    CCU2D add_134_29 (.A0(\register[2] [27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25812), .COUT(n25813), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_29.INIT0 = 16'h5aaa;
    defparam add_134_29.INIT1 = 16'h5aaa;
    defparam add_134_29.INJECT1_0 = "NO";
    defparam add_134_29.INJECT1_1 = "NO";
    CCU2D add_134_27 (.A0(\register[2] [25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25811), .COUT(n25812), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_27.INIT0 = 16'h5aaa;
    defparam add_134_27.INIT1 = 16'h5aaa;
    defparam add_134_27.INJECT1_0 = "NO";
    defparam add_134_27.INJECT1_1 = "NO";
    CCU2D add_134_25 (.A0(\register[2] [23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25810), .COUT(n25811), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_25.INIT0 = 16'h5aaa;
    defparam add_134_25.INIT1 = 16'h5aaa;
    defparam add_134_25.INJECT1_0 = "NO";
    defparam add_134_25.INJECT1_1 = "NO";
    CCU2D add_134_23 (.A0(\register[2] [21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25809), .COUT(n25810), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_23.INIT0 = 16'h5aaa;
    defparam add_134_23.INIT1 = 16'h5aaa;
    defparam add_134_23.INJECT1_0 = "NO";
    defparam add_134_23.INJECT1_1 = "NO";
    CCU2D add_134_21 (.A0(\register[2] [19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25808), .COUT(n25809), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_21.INIT0 = 16'h5aaa;
    defparam add_134_21.INIT1 = 16'h5aaa;
    defparam add_134_21.INJECT1_0 = "NO";
    defparam add_134_21.INJECT1_1 = "NO";
    LUT4 i21446_4_lut (.A(n30394), .B(\register_addr[2] ), .C(\register_addr[4] ), 
         .D(n9118), .Z(n28599)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21446_4_lut.init = 16'hfffe;
    CCU2D add_134_19 (.A0(\register[2] [17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25807), .COUT(n25808), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_19.INIT0 = 16'h5aaa;
    defparam add_134_19.INIT1 = 16'h5aaa;
    defparam add_134_19.INJECT1_0 = "NO";
    defparam add_134_19.INJECT1_1 = "NO";
    CCU2D add_134_17 (.A0(\register[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25806), .COUT(n25807), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_17.INIT0 = 16'h5aaa;
    defparam add_134_17.INIT1 = 16'h5aaa;
    defparam add_134_17.INJECT1_0 = "NO";
    defparam add_134_17.INJECT1_1 = "NO";
    CCU2D add_134_15 (.A0(\register[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25805), .COUT(n25806), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_15.INIT0 = 16'h5aaa;
    defparam add_134_15.INIT1 = 16'h5aaa;
    defparam add_134_15.INJECT1_0 = "NO";
    defparam add_134_15.INJECT1_1 = "NO";
    CCU2D add_134_13 (.A0(\register[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25804), .COUT(n25805), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_13.INIT0 = 16'h5aaa;
    defparam add_134_13.INIT1 = 16'h5aaa;
    defparam add_134_13.INJECT1_0 = "NO";
    defparam add_134_13.INJECT1_1 = "NO";
    CCU2D add_134_11 (.A0(\register[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25803), .COUT(n25804), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_11.INIT0 = 16'h5aaa;
    defparam add_134_11.INIT1 = 16'h5aaa;
    defparam add_134_11.INJECT1_0 = "NO";
    defparam add_134_11.INJECT1_1 = "NO";
    CCU2D add_134_9 (.A0(\register[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25802), .COUT(n25803), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_9.INIT0 = 16'h5aaa;
    defparam add_134_9.INIT1 = 16'h5aaa;
    defparam add_134_9.INJECT1_0 = "NO";
    defparam add_134_9.INJECT1_1 = "NO";
    CCU2D add_134_7 (.A0(\register[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25801), .COUT(n25802), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_7.INIT0 = 16'h5aaa;
    defparam add_134_7.INIT1 = 16'h5aaa;
    defparam add_134_7.INJECT1_0 = "NO";
    defparam add_134_7.INJECT1_1 = "NO";
    LUT4 i14633_3_lut (.A(\register[2] [3]), .B(n26507), .C(n30330), .Z(n5772[3])) /* synthesis lut_function=(!(A (B (C))+!A (B))) */ ;
    defparam i14633_3_lut.init = 16'h3b3b;
    CCU2D add_134_5 (.A0(\register[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25800), .COUT(n25801), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_5.INIT0 = 16'h5aaa;
    defparam add_134_5.INIT1 = 16'h5aaa;
    defparam add_134_5.INJECT1_0 = "NO";
    defparam add_134_5.INJECT1_1 = "NO";
    CCU2D add_134_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25799), .COUT(n25800), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_3.INIT0 = 16'h5aaa;
    defparam add_134_3.INIT1 = 16'h5aaa;
    defparam add_134_3.INJECT1_0 = "NO";
    defparam add_134_3.INJECT1_1 = "NO";
    CCU2D add_134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25799), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_1.INIT0 = 16'hF000;
    defparam add_134_1.INIT1 = 16'h5555;
    defparam add_134_1.INJECT1_0 = "NO";
    defparam add_134_1.INJECT1_1 = "NO";
    LUT4 i14778_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [5]), 
         .Z(n5772[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14778_2_lut_3_lut.init = 16'h2020;
    FD1P3IX read_size_i0_i1 (.D(n26670), .SP(n30307), .CD(n16116), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n30366), .SP(n30307), .CD(n16115), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    LUT4 i14792_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [4]), 
         .Z(n5772[4])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14792_2_lut_3_lut.init = 16'h2020;
    LUT4 i14549_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [14]), 
         .Z(n5772[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14549_2_lut_3_lut.init = 16'h2020;
    LUT4 i14581_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [17]), 
         .Z(n5772[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14581_2_lut_3_lut.init = 16'h2020;
    LUT4 i14553_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [12]), 
         .Z(n5772[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14553_2_lut_3_lut.init = 16'h2020;
    LUT4 i14557_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [10]), 
         .Z(n5772[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14557_2_lut_3_lut.init = 16'h2020;
    LUT4 i14401_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [8]), 
         .Z(n5772[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14401_2_lut_3_lut.init = 16'h2020;
    LUT4 i14504_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [16]), 
         .Z(n5772[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14504_2_lut_3_lut.init = 16'h2020;
    FD1P3AX read_value__i1 (.D(n29650), .SP(n30307), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3AX read_value__i2 (.D(n29613), .SP(n30307), .CK(debug_c_c), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5772[3]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5772[4]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n5772[5]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n5772[6]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n5772[7]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n5772[8]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n5772[9]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n5772[10]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n5772[11]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n5772[12]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n5772[13]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n5772[14]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n5772[15]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n5772[16]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n5772[17]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n5772[18]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n5772[19]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n5772[20]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n5772[21]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n5772[22]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n5772[23]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n5772[24]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n5772[25]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n5772[26]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n5772[27]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n5772[28]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n5772[29]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n5772[30]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n5772[31]), .SP(n30307), .CD(n9118), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_457 (.A(n28218), .B(n30324), .C(\register_addr[5] ), 
         .D(n30489), .Z(n8890)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(64[8] 95[15])
    defparam i2_4_lut_adj_457.init = 16'h0008;
    LUT4 i14554_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [11]), 
         .Z(n5772[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14554_2_lut_3_lut.init = 16'h2020;
    LUT4 i15029_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [20]), 
         .Z(n5772[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15029_2_lut_3_lut.init = 16'h2020;
    LUT4 i14791_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [6]), 
         .Z(n5772[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14791_2_lut_3_lut.init = 16'h2020;
    LUT4 i15122_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [18]), 
         .Z(n5772[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15122_2_lut_3_lut.init = 16'h2020;
    LUT4 i15033_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [19]), 
         .Z(n5772[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15033_2_lut_3_lut.init = 16'h2020;
    LUT4 i14550_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [13]), 
         .Z(n5772[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14550_2_lut_3_lut.init = 16'h2020;
    LUT4 i14495_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [9]), 
         .Z(n5772[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i14495_2_lut_3_lut.init = 16'h2020;
    LUT4 n29612_bdd_2_lut (.A(n29612), .B(n28599), .Z(n29613)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n29612_bdd_2_lut.init = 16'h2222;
    LUT4 register_addr_0__bdd_4_lut_22057 (.A(\register_addr[0] ), .B(\register[0] [2]), 
         .C(\register_addr[1] ), .D(\register[2] [2]), .Z(n29612)) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam register_addr_0__bdd_4_lut_22057.init = 16'h5e0e;
    LUT4 n29649_bdd_2_lut (.A(n29649), .B(n28599), .Z(n29650)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n29649_bdd_2_lut.init = 16'h2222;
    LUT4 i15025_2_lut_3_lut (.A(n26507), .B(n30330), .C(\register[2] [21]), 
         .Z(n5772[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15025_2_lut_3_lut.init = 16'h2020;
    \ClockDividerP(factor=12000000)  uptime_div (.clk_1Hz(clk_1Hz), .debug_c_c(debug_c_c), 
            .n32385(n32385), .GND_net(GND_net), .n32380(n32380)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(107[28] 109[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (clk_1Hz, debug_c_c, n32385, GND_net, 
            n32380) /* synthesis syn_module_defined=1 */ ;
    output clk_1Hz;
    input debug_c_c;
    input n32385;
    input GND_net;
    input n32380;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7608;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n2686;
    wire [31:0]n134;
    
    wire n26273, n26272, n26271, n26270, n26269, n26268, n26267, 
        n26266, n26265, n28706, n27, n26452, n25, n26, n24, 
        n19, n32, n28, n20, n26264, n26263, n26262, n29, n26_adj_516, 
        n26070, n26069, n26068, n26067, n26066, n26065, n26064, 
        n26063, n26062, n26061, n26060, n26059, n26058, n26057, 
        n26056, n26055;
    
    FD1S3IX clk_o_14 (.D(n7608), .CK(debug_c_c), .CD(n32385), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2610__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2686), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i0.GSR = "ENABLED";
    CCU2D add_19121_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26273), 
          .S0(n7608));
    defparam add_19121_cout.INIT0 = 16'h0000;
    defparam add_19121_cout.INIT1 = 16'h0000;
    defparam add_19121_cout.INJECT1_0 = "NO";
    defparam add_19121_cout.INJECT1_1 = "NO";
    CCU2D add_19121_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26272), .COUT(n26273));
    defparam add_19121_24.INIT0 = 16'h5555;
    defparam add_19121_24.INIT1 = 16'h5555;
    defparam add_19121_24.INJECT1_0 = "NO";
    defparam add_19121_24.INJECT1_1 = "NO";
    FD1S3IX count_2610__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2686), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i1.GSR = "ENABLED";
    CCU2D add_19121_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26271), .COUT(n26272));
    defparam add_19121_22.INIT0 = 16'h5555;
    defparam add_19121_22.INIT1 = 16'h5555;
    defparam add_19121_22.INJECT1_0 = "NO";
    defparam add_19121_22.INJECT1_1 = "NO";
    CCU2D add_19121_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26270), .COUT(n26271));
    defparam add_19121_20.INIT0 = 16'h5555;
    defparam add_19121_20.INIT1 = 16'h5555;
    defparam add_19121_20.INJECT1_0 = "NO";
    defparam add_19121_20.INJECT1_1 = "NO";
    CCU2D add_19121_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26269), .COUT(n26270));
    defparam add_19121_18.INIT0 = 16'h5555;
    defparam add_19121_18.INIT1 = 16'h5555;
    defparam add_19121_18.INJECT1_0 = "NO";
    defparam add_19121_18.INJECT1_1 = "NO";
    CCU2D add_19121_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26268), .COUT(n26269));
    defparam add_19121_16.INIT0 = 16'h5aaa;
    defparam add_19121_16.INIT1 = 16'h5555;
    defparam add_19121_16.INJECT1_0 = "NO";
    defparam add_19121_16.INJECT1_1 = "NO";
    CCU2D add_19121_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26267), .COUT(n26268));
    defparam add_19121_14.INIT0 = 16'h5aaa;
    defparam add_19121_14.INIT1 = 16'h5555;
    defparam add_19121_14.INJECT1_0 = "NO";
    defparam add_19121_14.INJECT1_1 = "NO";
    CCU2D add_19121_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26266), .COUT(n26267));
    defparam add_19121_12.INIT0 = 16'h5555;
    defparam add_19121_12.INIT1 = 16'h5aaa;
    defparam add_19121_12.INJECT1_0 = "NO";
    defparam add_19121_12.INJECT1_1 = "NO";
    CCU2D add_19121_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26265), .COUT(n26266));
    defparam add_19121_10.INIT0 = 16'h5aaa;
    defparam add_19121_10.INIT1 = 16'h5aaa;
    defparam add_19121_10.INJECT1_0 = "NO";
    defparam add_19121_10.INJECT1_1 = "NO";
    LUT4 i21656_2_lut (.A(n28706), .B(n32380), .Z(n2686)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21656_2_lut.init = 16'heeee;
    LUT4 i21654_4_lut (.A(n27), .B(n26452), .C(n25), .D(n26), .Z(n28706)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i21654_4_lut.init = 16'h0004;
    FD1S3IX count_2610__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2686), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i2.GSR = "ENABLED";
    FD1S3IX count_2610__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2686), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i3.GSR = "ENABLED";
    FD1S3IX count_2610__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2686), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i4.GSR = "ENABLED";
    FD1S3IX count_2610__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2686), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i5.GSR = "ENABLED";
    FD1S3IX count_2610__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2686), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i6.GSR = "ENABLED";
    FD1S3IX count_2610__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2686), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i7.GSR = "ENABLED";
    FD1S3IX count_2610__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2686), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i8.GSR = "ENABLED";
    FD1S3IX count_2610__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2686), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i9.GSR = "ENABLED";
    FD1S3IX count_2610__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i10.GSR = "ENABLED";
    FD1S3IX count_2610__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i11.GSR = "ENABLED";
    FD1S3IX count_2610__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i12.GSR = "ENABLED";
    FD1S3IX count_2610__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i13.GSR = "ENABLED";
    FD1S3IX count_2610__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i14.GSR = "ENABLED";
    FD1S3IX count_2610__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i15.GSR = "ENABLED";
    FD1S3IX count_2610__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i16.GSR = "ENABLED";
    FD1S3IX count_2610__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i17.GSR = "ENABLED";
    FD1S3IX count_2610__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i18.GSR = "ENABLED";
    FD1S3IX count_2610__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i19.GSR = "ENABLED";
    FD1S3IX count_2610__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i20.GSR = "ENABLED";
    FD1S3IX count_2610__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i21.GSR = "ENABLED";
    FD1S3IX count_2610__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i22.GSR = "ENABLED";
    FD1S3IX count_2610__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i23.GSR = "ENABLED";
    FD1S3IX count_2610__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i24.GSR = "ENABLED";
    FD1S3IX count_2610__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i25.GSR = "ENABLED";
    FD1S3IX count_2610__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i26.GSR = "ENABLED";
    FD1S3IX count_2610__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i27.GSR = "ENABLED";
    FD1S3IX count_2610__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i28.GSR = "ENABLED";
    FD1S3IX count_2610__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i29.GSR = "ENABLED";
    FD1S3IX count_2610__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i30.GSR = "ENABLED";
    FD1S3IX count_2610__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2686), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610__i31.GSR = "ENABLED";
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n26452)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    CCU2D add_19121_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26264), .COUT(n26265));
    defparam add_19121_8.INIT0 = 16'h5555;
    defparam add_19121_8.INIT1 = 16'h5aaa;
    defparam add_19121_8.INJECT1_0 = "NO";
    defparam add_19121_8.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    CCU2D add_19121_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26263), .COUT(n26264));
    defparam add_19121_6.INIT0 = 16'h5555;
    defparam add_19121_6.INIT1 = 16'h5555;
    defparam add_19121_6.INJECT1_0 = "NO";
    defparam add_19121_6.INJECT1_1 = "NO";
    CCU2D add_19121_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26262), .COUT(n26263));
    defparam add_19121_4.INIT0 = 16'h5aaa;
    defparam add_19121_4.INIT1 = 16'h5aaa;
    defparam add_19121_4.INJECT1_0 = "NO";
    defparam add_19121_4.INJECT1_1 = "NO";
    CCU2D add_19121_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26262));
    defparam add_19121_2.INIT0 = 16'h7000;
    defparam add_19121_2.INIT1 = 16'h5555;
    defparam add_19121_2.INJECT1_0 = "NO";
    defparam add_19121_2.INJECT1_1 = "NO";
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_516), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_451 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_451.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_452 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_452.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_516)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    CCU2D count_2610_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26070), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_33.INIT1 = 16'h0000;
    defparam count_2610_add_4_33.INJECT1_0 = "NO";
    defparam count_2610_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26069), .COUT(n26070), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_31.INJECT1_0 = "NO";
    defparam count_2610_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26068), .COUT(n26069), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_29.INJECT1_0 = "NO";
    defparam count_2610_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26067), .COUT(n26068), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_27.INJECT1_0 = "NO";
    defparam count_2610_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26066), .COUT(n26067), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_25.INJECT1_0 = "NO";
    defparam count_2610_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26065), .COUT(n26066), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_23.INJECT1_0 = "NO";
    defparam count_2610_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26064), .COUT(n26065), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_21.INJECT1_0 = "NO";
    defparam count_2610_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26063), .COUT(n26064), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_19.INJECT1_0 = "NO";
    defparam count_2610_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26062), .COUT(n26063), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_17.INJECT1_0 = "NO";
    defparam count_2610_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26061), .COUT(n26062), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_15.INJECT1_0 = "NO";
    defparam count_2610_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26060), .COUT(n26061), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_13.INJECT1_0 = "NO";
    defparam count_2610_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26059), .COUT(n26060), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_11.INJECT1_0 = "NO";
    defparam count_2610_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26058), .COUT(n26059), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_9.INJECT1_0 = "NO";
    defparam count_2610_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26057), .COUT(n26058), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_7.INJECT1_0 = "NO";
    defparam count_2610_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26056), .COUT(n26057), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_5.INJECT1_0 = "NO";
    defparam count_2610_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26055), .COUT(n26056), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2610_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2610_add_4_3.INJECT1_0 = "NO";
    defparam count_2610_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2610_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26055), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2610_add_4_1.INIT0 = 16'hF000;
    defparam count_2610_add_4_1.INIT1 = 16'h0555;
    defparam count_2610_add_4_1.INJECT1_0 = "NO";
    defparam count_2610_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module EncoderPeripheral_U11
//

module EncoderPeripheral_U11 (prev_select, debug_c_c, n30358, \register_addr[0] , 
            n30340, n30406, n30422, n30445, rw, n30349, n32380, 
            n9122, \quadA_delayed[1] , qreset, n6, \quadB_delayed[1] , 
            n14013, debug_c_0, encoder_li_c, encoder_lb_c, encoder_la_c, 
            \read_size[2] , n14291, n30366, read_value, \read_size[0] , 
            n302, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output prev_select;
    input debug_c_c;
    input n30358;
    input \register_addr[0] ;
    input n30340;
    input n30406;
    input n30422;
    input n30445;
    input rw;
    output n30349;
    input n32380;
    output n9122;
    input \quadA_delayed[1] ;
    output qreset;
    input n6;
    input \quadB_delayed[1] ;
    output n14013;
    input debug_c_0;
    input encoder_li_c;
    input encoder_lb_c;
    input encoder_la_c;
    output \read_size[2] ;
    input n14291;
    input n30366;
    output [31:0]read_value;
    output \read_size[0] ;
    input n302;
    input GND_net;
    input VCC_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    wire n28124, n28130, n28123, n28120, n28111, n28115, n28133, 
        n28112, n28125, n28126, n28128, n28129, n28127, n28121, 
        n28109, n28119, n28108, n28118, n28107, n28117, n28113, 
        n28122, n28110, n28116, n28114, n28106, n28132, n28131, 
        n28105;
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n6_adj_514;
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n14536;
    wire [31:0]n180;
    
    FD1S3AX prev_select_126 (.D(n30358), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam prev_select_126.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [4]), 
         .Z(n28124)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_422 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [5]), 
         .Z(n28130)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_422.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_423 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [6]), 
         .Z(n28123)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_423.init = 16'h2020;
    LUT4 i2_3_lut_rep_340_4_lut (.A(n30406), .B(n30422), .C(n30445), .D(rw), 
         .Z(n30349)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(78[9:33])
    defparam i2_3_lut_rep_340_4_lut.init = 16'h0010;
    LUT4 i2_3_lut_3_lut_4_lut (.A(n30406), .B(n30422), .C(n30445), .D(n32380), 
         .Z(n9122)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(78[9:33])
    defparam i2_3_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut_3_lut_adj_424 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [7]), 
         .Z(n28120)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_424.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_425 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [8]), 
         .Z(n28111)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_425.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_426 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [9]), 
         .Z(n28115)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_426.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_427 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [10]), 
         .Z(n28133)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_427.init = 16'h2020;
    LUT4 i1_4_lut (.A(\quadA_delayed[1] ), .B(qreset), .C(n6), .D(\quadB_delayed[1] ), 
         .Z(n14013)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(63[18:35])
    defparam i1_4_lut.init = 16'hedde;
    LUT4 i1_2_lut_3_lut_adj_428 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [11]), 
         .Z(n28112)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_428.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_429 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [12]), 
         .Z(n28125)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_429.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_430 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [13]), 
         .Z(n28126)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_430.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_431 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [14]), 
         .Z(n28128)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_431.init = 16'h2020;
    LUT4 i1_2_lut (.A(n32380), .B(debug_c_0), .Z(qreset)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(63[18:35])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_432 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [15]), 
         .Z(n28129)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_432.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_433 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [16]), 
         .Z(n28127)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_433.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_434 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [17]), 
         .Z(n28121)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_434.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_435 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [18]), 
         .Z(n28109)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_435.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_436 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [19]), 
         .Z(n28119)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_436.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_437 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [20]), 
         .Z(n28108)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_437.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_438 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [21]), 
         .Z(n28118)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_438.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_439 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [22]), 
         .Z(n28107)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_439.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_440 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [23]), 
         .Z(n28117)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_440.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_441 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [24]), 
         .Z(n28113)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_441.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_442 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [25]), 
         .Z(n28122)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_442.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_443 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [26]), 
         .Z(n28110)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_443.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_444 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [27]), 
         .Z(n28116)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_444.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_445 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [28]), 
         .Z(n28114)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_445.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_446 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [29]), 
         .Z(n28106)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_446.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_447 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [30]), 
         .Z(n28132)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_447.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_448 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [31]), 
         .Z(n28131)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_448.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_449 (.A(\register_addr[0] ), .B(n30340), .C(\register[1] [0]), 
         .Z(n28105)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_449.init = 16'h2020;
    LUT4 i1_4_lut_adj_450 (.A(quadA_delayed[1]), .B(qreset), .C(n6_adj_514), 
         .D(quadB_delayed[1]), .Z(n14536)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(63[18:35])
    defparam i1_4_lut_adj_450.init = 16'hedde;
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_li_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n180[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_lb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n180[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_la_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n180[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_size__i2 (.D(n30366), .SP(n14291), .CD(n30340), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n180[1]), .SP(n14291), .CD(n30340), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n180[2]), .SP(n14291), .CD(n30340), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n180[3]), .SP(n14291), .CD(n30340), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n28124), .SP(n14291), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n28130), .SP(n14291), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n28123), .SP(n14291), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n28120), .SP(n14291), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n28111), .SP(n14291), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n28115), .SP(n14291), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n28133), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n28112), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n28125), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n28126), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n28128), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n28129), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n28127), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n28121), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n28109), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n28119), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n28108), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n28118), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n28107), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n28117), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n28113), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n28122), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n28110), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n28116), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n28114), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n28106), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n28132), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n28131), .SP(n14291), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_size__i1 (.D(n302), .SP(n14291), .CD(n30340), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX read_value__i0 (.D(n28105), .SP(n14291), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=649, LSE_RLINE=659 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i0.GSR = "ENABLED";
    QuadratureDecoder_U6 q (.quadA_delayed({Open_7, quadA_delayed[1], Open_8}), 
            .GND_net(GND_net), .n6(n6_adj_514), .\register[1] ({\register[1] }), 
            .debug_c_c(debug_c_c), .qreset(qreset), .VCC_net(VCC_net), 
            .encoder_lb_c(encoder_lb_c), .encoder_la_c(encoder_la_c), .n14536(n14536), 
            .\quadB_delayed[1] (quadB_delayed[1])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(93[20] 97[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder_U6
//

module QuadratureDecoder_U6 (quadA_delayed, GND_net, n6, \register[1] , 
            debug_c_c, qreset, VCC_net, encoder_lb_c, encoder_la_c, 
            n14536, \quadB_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    output [2:0]quadA_delayed;
    input GND_net;
    output n6;
    output [31:0]\register[1] ;
    input debug_c_c;
    input qreset;
    input VCC_net;
    input encoder_lb_c;
    input encoder_la_c;
    input n14536;
    output \quadB_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25605;
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [31:0]n100;
    
    wire n25604, n25603, n25602, n25601, n25600, n25599;
    wire [2:0]quadA_delayed_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n25598, n25597, n25596, n25595, n25594, n25593, n25592, 
        n25591, n25590;
    wire [31:0]n4222;
    
    CCU2D add_1683_33 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n25605), .S0(n100[30]), 
          .S1(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_33.INIT0 = 16'h6969;
    defparam add_1683_33.INIT1 = 16'h6969;
    defparam add_1683_33.INJECT1_0 = "NO";
    defparam add_1683_33.INJECT1_1 = "NO";
    CCU2D add_1683_31 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n25604), .COUT(n25605), 
          .S0(n100[28]), .S1(n100[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_31.INIT0 = 16'h6969;
    defparam add_1683_31.INIT1 = 16'h6969;
    defparam add_1683_31.INJECT1_0 = "NO";
    defparam add_1683_31.INJECT1_1 = "NO";
    CCU2D add_1683_29 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n25603), .COUT(n25604), 
          .S0(n100[26]), .S1(n100[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_29.INIT0 = 16'h6969;
    defparam add_1683_29.INIT1 = 16'h6969;
    defparam add_1683_29.INJECT1_0 = "NO";
    defparam add_1683_29.INJECT1_1 = "NO";
    CCU2D add_1683_27 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n25602), .COUT(n25603), 
          .S0(n100[24]), .S1(n100[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_27.INIT0 = 16'h6969;
    defparam add_1683_27.INIT1 = 16'h6969;
    defparam add_1683_27.INJECT1_0 = "NO";
    defparam add_1683_27.INJECT1_1 = "NO";
    CCU2D add_1683_25 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n25601), .COUT(n25602), 
          .S0(n100[22]), .S1(n100[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_25.INIT0 = 16'h6969;
    defparam add_1683_25.INIT1 = 16'h6969;
    defparam add_1683_25.INJECT1_0 = "NO";
    defparam add_1683_25.INJECT1_1 = "NO";
    CCU2D add_1683_23 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n25600), .COUT(n25601), 
          .S0(n100[20]), .S1(n100[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_23.INIT0 = 16'h6969;
    defparam add_1683_23.INIT1 = 16'h6969;
    defparam add_1683_23.INJECT1_0 = "NO";
    defparam add_1683_23.INJECT1_1 = "NO";
    CCU2D add_1683_21 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n25599), .COUT(n25600), 
          .S0(n100[18]), .S1(n100[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_21.INIT0 = 16'h6969;
    defparam add_1683_21.INIT1 = 16'h6969;
    defparam add_1683_21.INJECT1_0 = "NO";
    defparam add_1683_21.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed_c[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    CCU2D add_1683_19 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n25598), .COUT(n25599), 
          .S0(n100[16]), .S1(n100[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_19.INIT0 = 16'h6969;
    defparam add_1683_19.INIT1 = 16'h6969;
    defparam add_1683_19.INJECT1_0 = "NO";
    defparam add_1683_19.INJECT1_1 = "NO";
    CCU2D add_1683_17 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n25597), .COUT(n25598), 
          .S0(n100[14]), .S1(n100[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_17.INIT0 = 16'h6969;
    defparam add_1683_17.INIT1 = 16'h6969;
    defparam add_1683_17.INJECT1_0 = "NO";
    defparam add_1683_17.INJECT1_1 = "NO";
    CCU2D add_1683_15 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n25596), .COUT(n25597), 
          .S0(n100[12]), .S1(n100[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_15.INIT0 = 16'h6969;
    defparam add_1683_15.INIT1 = 16'h6969;
    defparam add_1683_15.INJECT1_0 = "NO";
    defparam add_1683_15.INJECT1_1 = "NO";
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_lb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_la_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed_c[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    CCU2D add_1683_13 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n25595), .COUT(n25596), 
          .S0(n100[10]), .S1(n100[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_13.INIT0 = 16'h6969;
    defparam add_1683_13.INIT1 = 16'h6969;
    defparam add_1683_13.INJECT1_0 = "NO";
    defparam add_1683_13.INJECT1_1 = "NO";
    CCU2D add_1683_11 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n25594), .COUT(n25595), 
          .S0(n100[8]), .S1(n100[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_11.INIT0 = 16'h6969;
    defparam add_1683_11.INIT1 = 16'h6969;
    defparam add_1683_11.INJECT1_0 = "NO";
    defparam add_1683_11.INJECT1_1 = "NO";
    CCU2D add_1683_9 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n25593), .COUT(n25594), 
          .S0(n100[6]), .S1(n100[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_9.INIT0 = 16'h6969;
    defparam add_1683_9.INIT1 = 16'h6969;
    defparam add_1683_9.INJECT1_0 = "NO";
    defparam add_1683_9.INJECT1_1 = "NO";
    CCU2D add_1683_7 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n25592), .COUT(n25593), 
          .S0(n100[4]), .S1(n100[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_7.INIT0 = 16'h6969;
    defparam add_1683_7.INIT1 = 16'h6969;
    defparam add_1683_7.INJECT1_0 = "NO";
    defparam add_1683_7.INJECT1_1 = "NO";
    CCU2D add_1683_5 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n25591), .COUT(n25592), 
          .S0(n100[2]), .S1(n100[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_5.INIT0 = 16'h6969;
    defparam add_1683_5.INIT1 = 16'h6969;
    defparam add_1683_5.INJECT1_0 = "NO";
    defparam add_1683_5.INJECT1_1 = "NO";
    CCU2D add_1683_3 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n25590), .COUT(n25591), 
          .S0(n4222[0]), .S1(n4222[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_3.INIT0 = 16'h9696;
    defparam add_1683_3.INIT1 = 16'h6969;
    defparam add_1683_3.INJECT1_0 = "NO";
    defparam add_1683_3.INJECT1_1 = "NO";
    CCU2D add_1683_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n25590));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1683_1.INIT0 = 16'hF000;
    defparam add_1683_1.INIT1 = 16'h6666;
    defparam add_1683_1.INJECT1_0 = "NO";
    defparam add_1683_1.INJECT1_1 = "NO";
    FD1P3IX count__i1 (.D(n4222[1]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i0 (.D(n4222[0]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n100[2]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n100[3]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n100[4]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n100[5]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n100[6]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n100[7]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n100[8]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n100[9]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n100[10]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n100[11]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n100[12]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n100[13]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n100[14]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n100[15]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n100[16]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n100[17]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n100[18]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n100[19]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n100[20]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n100[21]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n100[22]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n100[23]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n100[24]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n100[25]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n100[26]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n100[27]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n100[28]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n100[29]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n100[30]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i31 (.D(n100[31]), .SP(n14536), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed_c[0]), .CK(debug_c_c), .Q(quadA_delayed[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(quadA_delayed[1]), .CK(debug_c_c), .Q(quadA_delayed_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP_SP(factor=120000) 
//

module \ClockDividerP_SP(factor=120000)  (GND_net, debug_c_0, debug_c_c, 
            n32385, n32380) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output debug_c_0;
    input debug_c_c;
    input n32385;
    input n32380;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30356, n20, n19, n21, n26840, n26038;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(86[13:18])
    wire [31:0]n134;
    
    wire n26037, n26036, n26035, n26034, n26033, n26032, n26031, 
        n26030, n26029, n26028, n26027, n26026, n26025, n26024, 
        n26023, n2676, n25, n38, n34, n26, n28709, n28413, n28595, 
        n28411, n28569, n28419, n36, n30, n32, n22;
    
    LUT4 i21727_4_lut_4_lut (.A(n30356), .B(n20), .C(n19), .D(n21), 
         .Z(n26840)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i21727_4_lut_4_lut.init = 16'h0001;
    CCU2D count_2609_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26038), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_33.INIT1 = 16'h0000;
    defparam count_2609_add_4_33.INJECT1_0 = "NO";
    defparam count_2609_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26037), .COUT(n26038), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_31.INJECT1_0 = "NO";
    defparam count_2609_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26036), .COUT(n26037), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_29.INJECT1_0 = "NO";
    defparam count_2609_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26035), .COUT(n26036), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_27.INJECT1_0 = "NO";
    defparam count_2609_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26034), .COUT(n26035), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_25.INJECT1_0 = "NO";
    defparam count_2609_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26033), .COUT(n26034), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_23.INJECT1_0 = "NO";
    defparam count_2609_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26032), .COUT(n26033), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_21.INJECT1_0 = "NO";
    defparam count_2609_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26031), .COUT(n26032), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_19.INJECT1_0 = "NO";
    defparam count_2609_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26030), .COUT(n26031), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_17.INJECT1_0 = "NO";
    defparam count_2609_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26029), .COUT(n26030), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_15.INJECT1_0 = "NO";
    defparam count_2609_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26028), .COUT(n26029), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_13.INJECT1_0 = "NO";
    defparam count_2609_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26027), .COUT(n26028), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_11.INJECT1_0 = "NO";
    defparam count_2609_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26026), .COUT(n26027), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_9.INJECT1_0 = "NO";
    defparam count_2609_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26025), .COUT(n26026), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_7.INJECT1_0 = "NO";
    defparam count_2609_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26024), .COUT(n26025), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_5.INJECT1_0 = "NO";
    defparam count_2609_add_4_5.INJECT1_1 = "NO";
    FD1S3IX clk_o_13 (.D(n26840), .CK(debug_c_c), .CD(n32385), .Q(debug_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(88[9] 107[6])
    defparam clk_o_13.GSR = "ENABLED";
    CCU2D count_2609_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26023), .COUT(n26024), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2609_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2609_add_4_3.INJECT1_0 = "NO";
    defparam count_2609_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2609_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26023), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609_add_4_1.INIT0 = 16'hF000;
    defparam count_2609_add_4_1.INIT1 = 16'h0555;
    defparam count_2609_add_4_1.INJECT1_0 = "NO";
    defparam count_2609_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2609__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2676), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i0.GSR = "ENABLED";
    LUT4 i19_4_lut_rep_347 (.A(n25), .B(n38), .C(n34), .D(n26), .Z(n30356)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i19_4_lut_rep_347.init = 16'hfffe;
    LUT4 i21659_2_lut (.A(n28709), .B(n32380), .Z(n2676)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21659_2_lut.init = 16'heeee;
    LUT4 i21657_4_lut (.A(n30356), .B(n28413), .C(n28595), .D(n28411), 
         .Z(n28709)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i21657_4_lut.init = 16'h4000;
    LUT4 i21266_2_lut (.A(count[10]), .B(count[12]), .Z(n28413)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21266_2_lut.init = 16'h8888;
    LUT4 i21442_4_lut (.A(count[3]), .B(n28569), .C(n28419), .D(count[0]), 
         .Z(n28595)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i21442_4_lut.init = 16'h8000;
    LUT4 i21264_2_lut (.A(count[2]), .B(count[5]), .Z(n28411)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21264_2_lut.init = 16'h8888;
    LUT4 i21416_4_lut (.A(count[1]), .B(count[16]), .C(count[4]), .D(count[15]), 
         .Z(n28569)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i21416_4_lut.init = 16'h8000;
    LUT4 i21272_2_lut (.A(count[7]), .B(count[14]), .Z(n28419)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21272_2_lut.init = 16'h8888;
    FD1S3IX count_2609__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2676), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i1.GSR = "ENABLED";
    FD1S3IX count_2609__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2676), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i2.GSR = "ENABLED";
    FD1S3IX count_2609__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2676), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i3.GSR = "ENABLED";
    FD1S3IX count_2609__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2676), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i4.GSR = "ENABLED";
    FD1S3IX count_2609__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2676), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i5.GSR = "ENABLED";
    FD1S3IX count_2609__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2676), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i6.GSR = "ENABLED";
    FD1S3IX count_2609__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2676), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i7.GSR = "ENABLED";
    FD1S3IX count_2609__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2676), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i8.GSR = "ENABLED";
    FD1S3IX count_2609__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2676), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i9.GSR = "ENABLED";
    FD1S3IX count_2609__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i10.GSR = "ENABLED";
    FD1S3IX count_2609__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i11.GSR = "ENABLED";
    FD1S3IX count_2609__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i12.GSR = "ENABLED";
    FD1S3IX count_2609__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i13.GSR = "ENABLED";
    FD1S3IX count_2609__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i14.GSR = "ENABLED";
    FD1S3IX count_2609__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i15.GSR = "ENABLED";
    FD1S3IX count_2609__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i16.GSR = "ENABLED";
    FD1S3IX count_2609__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i17.GSR = "ENABLED";
    FD1S3IX count_2609__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i18.GSR = "ENABLED";
    FD1S3IX count_2609__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i19.GSR = "ENABLED";
    FD1S3IX count_2609__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i20.GSR = "ENABLED";
    FD1S3IX count_2609__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i21.GSR = "ENABLED";
    FD1S3IX count_2609__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i22.GSR = "ENABLED";
    FD1S3IX count_2609__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i23.GSR = "ENABLED";
    FD1S3IX count_2609__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i24.GSR = "ENABLED";
    FD1S3IX count_2609__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i25.GSR = "ENABLED";
    FD1S3IX count_2609__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i26.GSR = "ENABLED";
    FD1S3IX count_2609__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i27.GSR = "ENABLED";
    FD1S3IX count_2609__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i28.GSR = "ENABLED";
    FD1S3IX count_2609__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i29.GSR = "ENABLED";
    FD1S3IX count_2609__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i30.GSR = "ENABLED";
    FD1S3IX count_2609__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2676), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2609__i31.GSR = "ENABLED";
    LUT4 i9_4_lut (.A(count[5]), .B(count[16]), .C(count[12]), .D(count[14]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(count[7]), .B(count[15]), .C(count[4]), .D(count[10]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[1]), .B(count[0]), .C(count[2]), .D(count[3]), 
         .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[11]), .B(count[13]), .Z(n25)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(count[6]), .B(n36), .C(n30), .D(count[9]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(count[20]), .B(count[31]), .C(count[24]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(count[21]), .B(count[17]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i16_4_lut (.A(count[26]), .B(n32), .C(n22), .D(count[29]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(count[18]), .B(count[28]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(count[25]), .B(count[23]), .C(count[8]), .D(count[27]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[19]), .B(count[22]), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i2_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (\register_addr[1] , \register_addr[0] , 
            debug_c_c, VCC_net, GND_net, Stepper_Z_nFault_c, n32382, 
            \read_size[0] , n13918, n28323, Stepper_Z_M0_c_0, n579, 
            prev_step_clk, step_clk, n13594, prev_select, n30391, 
            Stepper_Z_M2_c_2, n32, n30422, \register_addr[2] , n26507, 
            \register_addr[3] , n32380, n26486, read_value, \steps_reg[5] , 
            \steps_reg[6] , \steps_reg[9] , \steps_reg[3] , databus, 
            n3892, n13269, \register_addr[4] , n30344, \register_addr[5] , 
            limit_c_2, n30421, int_step, n22, n30310, n30317, n32385, 
            n32381, n32386, \div_factor_reg[9] , \div_factor_reg[6] , 
            \div_factor_reg[5] , \div_factor_reg[3] , \control_reg[7] , 
            Stepper_Z_En_c, Stepper_Z_Dir_c, \control_reg[3] , Stepper_Z_M1_c_1, 
            \read_size[2] , n30342, n20670, n20681, n6917, n28148, 
            n8272) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[1] ;
    input \register_addr[0] ;
    input debug_c_c;
    input VCC_net;
    input GND_net;
    input Stepper_Z_nFault_c;
    input n32382;
    output \read_size[0] ;
    input n13918;
    input n28323;
    output Stepper_Z_M0_c_0;
    input n579;
    output prev_step_clk;
    output step_clk;
    input n13594;
    output prev_select;
    input n30391;
    output Stepper_Z_M2_c_2;
    input n32;
    input n30422;
    input \register_addr[2] ;
    output n26507;
    input \register_addr[3] ;
    input n32380;
    output n26486;
    output [31:0]read_value;
    output \steps_reg[5] ;
    output \steps_reg[6] ;
    output \steps_reg[9] ;
    output \steps_reg[3] ;
    input [31:0]databus;
    input n3892;
    input n13269;
    input \register_addr[4] ;
    input n30344;
    input \register_addr[5] ;
    input limit_c_2;
    input n30421;
    output int_step;
    input n22;
    input n30310;
    input n30317;
    input n32385;
    input n32381;
    input n32386;
    output \div_factor_reg[9] ;
    output \div_factor_reg[6] ;
    output \div_factor_reg[5] ;
    output \div_factor_reg[3] ;
    output \control_reg[7] ;
    output Stepper_Z_En_c;
    output Stepper_Z_Dir_c;
    output \control_reg[3] ;
    output Stepper_Z_M1_c_1;
    output \read_size[2] ;
    input n30342;
    input n20670;
    input n20681;
    input n6917;
    input n28148;
    input n8272;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n28155, n28156, fault_latched;
    wire [31:0]n3893;
    
    wire n21775, limit_latched, n182, prev_limit_latched, n28157, 
        n28158, n28640, n28641, n28642, n7, n11679, n49, n62, 
        n58, n50, n41, n60, n54, n42;
    wire [31:0]n100;
    
    wire n52, n38, n56, n46;
    wire [31:0]n224;
    
    wire n13591, n28171, n28150, n28151, n28152, n28153, n28159, 
        n28154, n28160, n28161, n28162, n28163, n28164, n28165, 
        n28166, n28167, n28673, n28674, n28675, n28168, n28149;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n28687;
    wire [31:0]n6891;
    
    wire n25934, n25933, n25932, n25931, n25930, n25929, n25928, 
        n25927, n25926, n25925, n25924, n25923, n25922, n25921, 
        n25920, n28685, n28686, n25919;
    wire [7:0]n8271;
    wire [31:0]n6855;
    
    LUT4 i1_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n28155)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_403 (.A(div_factor_reg[15]), .B(\register_addr[1] ), 
         .C(steps_reg[15]), .D(\register_addr[0] ), .Z(n28156)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_403.init = 16'hc088;
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3893[0]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n28323), .SP(n13918), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n21775), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13594), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n30391), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_404 (.A(div_factor_reg[16]), .B(\register_addr[1] ), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n28157)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_404.init = 16'hc088;
    LUT4 i1_4_lut_adj_405 (.A(div_factor_reg[20]), .B(\register_addr[1] ), 
         .C(steps_reg[20]), .D(\register_addr[0] ), .Z(n28158)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_405.init = 16'hc088;
    PFUMX i21489 (.BLUT(n28640), .ALUT(n28641), .C0(\register_addr[0] ), 
          .Z(n28642));
    LUT4 i21487_3_lut (.A(Stepper_Z_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n28640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21487_3_lut.init = 16'hcaca;
    LUT4 i21488_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n28641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21488_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut (.A(n7), .B(n30422), .C(\register_addr[2] ), .D(\register_addr[1] ), 
         .Z(n26507)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i4_4_lut.init = 16'hffef;
    LUT4 i2_2_lut (.A(\register_addr[3] ), .B(\register_addr[0] ), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i5272_3_lut (.A(prev_limit_latched), .B(n32380), .C(limit_latched), 
         .Z(n11679)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i5272_3_lut.init = 16'hdcdc;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n26486)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n13918), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n13918), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n13918), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1564_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3892), .Z(n3893[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i1_3_lut.init = 16'hcaca;
    LUT4 i21815_2_lut (.A(n13591), .B(n32380), .Z(n21775)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21815_2_lut.init = 16'heeee;
    LUT4 i21686_4_lut (.A(n13269), .B(\register_addr[4] ), .C(n30344), 
         .D(\register_addr[5] ), .Z(n13591)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i21686_4_lut.init = 16'h1000;
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n30421), .B(\register_addr[4] ), .C(\register_addr[5] ), 
         .Z(n28171)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i2_3_lut.init = 16'h2020;
    LUT4 mux_1564_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3892), 
         .Z(n3893[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3892), 
         .Z(n3893[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3892), 
         .Z(n3893[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3892), 
         .Z(n3893[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3892), 
         .Z(n3893[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3892), 
         .Z(n3893[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3892), 
         .Z(n3893[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3892), 
         .Z(n3893[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3892), 
         .Z(n3893[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3892), 
         .Z(n3893[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3892), 
         .Z(n3893[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3892), 
         .Z(n3893[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3892), 
         .Z(n3893[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3892), 
         .Z(n3893[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3892), 
         .Z(n3893[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3892), 
         .Z(n3893[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3892), 
         .Z(n3893[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3892), 
         .Z(n3893[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3892), 
         .Z(n3893[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3892), 
         .Z(n3893[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3892), 
         .Z(n3893[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3892), 
         .Z(n3893[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3892), .Z(n3893[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3892), .Z(n3893[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3892), .Z(n3893[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3892), .Z(n3893[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3892), .Z(n3893[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3892), .Z(n3893[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3892), .Z(n3893[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3892), .Z(n3893[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3892), .Z(n3893[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1564_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_406 (.A(div_factor_reg[8]), .B(\register_addr[1] ), 
         .C(steps_reg[8]), .D(\register_addr[0] ), .Z(n28150)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_406.init = 16'hc088;
    LUT4 i1_4_lut_adj_407 (.A(div_factor_reg[10]), .B(\register_addr[1] ), 
         .C(steps_reg[10]), .D(\register_addr[0] ), .Z(n28151)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_407.init = 16'hc088;
    LUT4 i1_4_lut_adj_408 (.A(div_factor_reg[11]), .B(\register_addr[1] ), 
         .C(steps_reg[11]), .D(\register_addr[0] ), .Z(n28152)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_408.init = 16'hc088;
    LUT4 i1_4_lut_adj_409 (.A(div_factor_reg[12]), .B(\register_addr[1] ), 
         .C(steps_reg[12]), .D(\register_addr[0] ), .Z(n28153)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_409.init = 16'hc088;
    LUT4 i1_4_lut_adj_410 (.A(div_factor_reg[21]), .B(\register_addr[1] ), 
         .C(steps_reg[21]), .D(\register_addr[0] ), .Z(n28159)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_410.init = 16'hc088;
    LUT4 i1_4_lut_adj_411 (.A(div_factor_reg[13]), .B(\register_addr[1] ), 
         .C(steps_reg[13]), .D(\register_addr[0] ), .Z(n28154)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_411.init = 16'hc088;
    LUT4 i1_4_lut_adj_412 (.A(div_factor_reg[22]), .B(\register_addr[1] ), 
         .C(steps_reg[22]), .D(\register_addr[0] ), .Z(n28160)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_412.init = 16'hc088;
    LUT4 i1_4_lut_adj_413 (.A(div_factor_reg[23]), .B(\register_addr[1] ), 
         .C(steps_reg[23]), .D(\register_addr[0] ), .Z(n28161)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_413.init = 16'hc088;
    LUT4 i1_4_lut_adj_414 (.A(div_factor_reg[24]), .B(\register_addr[1] ), 
         .C(steps_reg[24]), .D(\register_addr[0] ), .Z(n28162)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_414.init = 16'hc088;
    LUT4 i1_4_lut_adj_415 (.A(div_factor_reg[25]), .B(\register_addr[1] ), 
         .C(steps_reg[25]), .D(\register_addr[0] ), .Z(n28163)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_415.init = 16'hc088;
    LUT4 i1_4_lut_adj_416 (.A(div_factor_reg[26]), .B(\register_addr[1] ), 
         .C(steps_reg[26]), .D(\register_addr[0] ), .Z(n28164)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_416.init = 16'hc088;
    LUT4 i1_4_lut_adj_417 (.A(div_factor_reg[27]), .B(\register_addr[1] ), 
         .C(steps_reg[27]), .D(\register_addr[0] ), .Z(n28165)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_417.init = 16'hc088;
    FD1P3AX int_step_182 (.D(n30310), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_418 (.A(div_factor_reg[28]), .B(\register_addr[1] ), 
         .C(steps_reg[28]), .D(\register_addr[0] ), .Z(n28166)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_418.init = 16'hc088;
    LUT4 i1_4_lut_adj_419 (.A(div_factor_reg[29]), .B(\register_addr[1] ), 
         .C(steps_reg[29]), .D(\register_addr[0] ), .Z(n28167)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_419.init = 16'hc088;
    PFUMX i21522 (.BLUT(n28673), .ALUT(n28674), .C0(\register_addr[1] ), 
          .Z(n28675));
    LUT4 i1_4_lut_adj_420 (.A(div_factor_reg[30]), .B(\register_addr[1] ), 
         .C(steps_reg[30]), .D(\register_addr[0] ), .Z(n28168)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_420.init = 16'hc088;
    LUT4 i1_4_lut_adj_421 (.A(div_factor_reg[31]), .B(\register_addr[1] ), 
         .C(steps_reg[31]), .D(\register_addr[0] ), .Z(n28149)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_421.init = 16'hc088;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n30317), .CD(n32386), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n30317), .CD(n32386), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n30317), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n30317), .PD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n30317), .PD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n30317), .PD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n30317), .PD(n32381), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n30317), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n30317), .PD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n30317), .PD(n32385), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n30317), .PD(n32381), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n30317), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n30317), .CD(n32385), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13591), .CD(n11679), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13591), .PD(n32385), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13591), .PD(n32385), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13591), .CD(n32382), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13591), .PD(n32382), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13591), .CD(n32382), 
            .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13591), .PD(n32382), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n28171), .SP(n13918), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3893[31]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3893[30]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3893[29]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3893[28]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3893[27]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3893[26]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3893[25]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3893[24]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3893[23]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3893[22]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3893[21]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3893[20]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3893[19]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3893[18]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3893[17]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3893[16]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3893[15]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3893[14]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3893[13]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3893[12]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3893[11]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3893[10]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3893[9]), .CK(debug_c_c), .CD(n30342), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3893[8]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3893[7]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3893[6]), .CK(debug_c_c), .CD(n30342), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3893[5]), .CK(debug_c_c), .CD(n30342), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3893[4]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3893[3]), .CK(debug_c_c), .CD(n30342), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3893[2]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3893[1]), .CK(debug_c_c), .CD(n30342), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n28687), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i14614_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14614_4_lut.init = 16'hc088;
    LUT4 i14615_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14615_4_lut.init = 16'hc088;
    LUT4 i14616_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14616_4_lut.init = 16'hc088;
    FD1P3IX read_value__i2 (.D(n28642), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n20670), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6891[4]), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n20681), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6917), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6891[7]), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n28150), .SP(n13918), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n28148), .SP(n13918), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n28151), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n28152), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n28153), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n28154), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n28155), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n28156), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n28157), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n28158), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n28159), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n28160), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n28161), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n28162), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n28163), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n28164), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n28165), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n28166), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n28167), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n28168), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n28149), .SP(n13918), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25934), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25933), .COUT(n25934), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25932), .COUT(n25933), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25931), .COUT(n25932), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25930), .COUT(n25931), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25929), .COUT(n25930), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25928), .COUT(n25929), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25927), .COUT(n25928), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25926), .COUT(n25927), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25925), .COUT(n25926), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25924), .COUT(n25925), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25923), .COUT(n25924), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25922), .COUT(n25923), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25921), .COUT(n25922), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25920), .COUT(n25921), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 i21532_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n28685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21532_3_lut.init = 16'hcaca;
    LUT4 i21533_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n28686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21533_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25919), .COUT(n25920), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n25919), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    FD1P3IX read_value__i0 (.D(n28675), .SP(n13918), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i21520_3_lut (.A(Stepper_Z_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n28673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21520_3_lut.init = 16'hcaca;
    LUT4 i21521_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n28674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21521_3_lut.init = 16'hcaca;
    PFUMX i21534 (.BLUT(n28685), .ALUT(n28686), .C0(\register_addr[1] ), 
          .Z(n28687));
    LUT4 i14617_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8271[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14617_2_lut.init = 16'h2222;
    LUT4 mux_1941_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n6855[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1941_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1941_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6855[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1941_i8_3_lut.init = 16'hcaca;
    PFUMX mux_1945_i5 (.BLUT(n8271[4]), .ALUT(n6855[4]), .C0(\register_addr[1] ), 
          .Z(n6891[4]));
    PFUMX mux_1945_i8 (.BLUT(n8272), .ALUT(n6855[7]), .C0(\register_addr[1] ), 
          .Z(n6891[7]));
    ClockDivider step_clk_gen (.div_factor_reg({div_factor_reg[31:10], \div_factor_reg[9] , 
            div_factor_reg[8:7], \div_factor_reg[6] , \div_factor_reg[5] , 
            div_factor_reg[4], \div_factor_reg[3] , div_factor_reg[2:0]}), 
            .GND_net(GND_net), .n32380(n32380), .step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n32385(n32385)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (div_factor_reg, GND_net, n32380, step_clk, debug_c_c, 
            n32385) /* synthesis syn_module_defined=1 */ ;
    input [31:0]div_factor_reg;
    input GND_net;
    input n32380;
    output step_clk;
    input debug_c_c;
    input n32385;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25659, n25660, n25658, n7886, n30301, n7920, n16222, 
        n25657, n25656, n25655, n25870;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n25869, n7851, n25868, n26022;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n26021, n25867, n25866, n26020, n26019, n26018, n25865, 
        n25864, n26017, n26016, n25863, n26015, n25862, n26014, 
        n26013, n25861, n25860, n26012, n25859, n26011, n26010, 
        n26009, n25858, n26008, n26007, n25857, n25856, n25855, 
        n25702, n25701, n25700, n25699, n25698, n25697, n25696, 
        n25695, n25694, n25693, n25692, n25691, n25690, n25689, 
        n25688, n25687, n25686, n25685, n25684, n25683, n25682, 
        n25681, n25680, n25679, n25678, n25677, n25676, n25675, 
        n25674, n25673, n25672, n25671, n25670, n25669, n25668, 
        n25667, n25666, n25665, n25664, n25663, n25662, n25661;
    
    CCU2D sub_2027_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25659), .COUT(n25660));
    defparam sub_2027_add_2_11.INIT0 = 16'hf555;
    defparam sub_2027_add_2_11.INIT1 = 16'hf555;
    defparam sub_2027_add_2_11.INJECT1_0 = "NO";
    defparam sub_2027_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25658), .COUT(n25659));
    defparam sub_2027_add_2_9.INIT0 = 16'hf555;
    defparam sub_2027_add_2_9.INIT1 = 16'hf555;
    defparam sub_2027_add_2_9.INJECT1_0 = "NO";
    defparam sub_2027_add_2_9.INJECT1_1 = "NO";
    LUT4 i1017_2_lut_rep_292 (.A(n7886), .B(n32380), .Z(n30301)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1017_2_lut_rep_292.init = 16'heeee;
    LUT4 i9810_2_lut_3_lut (.A(n7886), .B(n32380), .C(n7920), .Z(n16222)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9810_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_2027_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25657), .COUT(n25658));
    defparam sub_2027_add_2_7.INIT0 = 16'hf555;
    defparam sub_2027_add_2_7.INIT1 = 16'hf555;
    defparam sub_2027_add_2_7.INJECT1_0 = "NO";
    defparam sub_2027_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25656), .COUT(n25657));
    defparam sub_2027_add_2_5.INIT0 = 16'hf555;
    defparam sub_2027_add_2_5.INIT1 = 16'hf555;
    defparam sub_2027_add_2_5.INJECT1_0 = "NO";
    defparam sub_2027_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25655), .COUT(n25656));
    defparam sub_2027_add_2_3.INIT0 = 16'hf555;
    defparam sub_2027_add_2_3.INIT1 = 16'hf555;
    defparam sub_2027_add_2_3.INJECT1_0 = "NO";
    defparam sub_2027_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n25655));
    defparam sub_2027_add_2_1.INIT0 = 16'h0000;
    defparam sub_2027_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2027_add_2_1.INJECT1_0 = "NO";
    defparam sub_2027_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25870), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25869), .COUT(n25870), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7851), .CK(debug_c_c), .CD(n32385), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25868), .COUT(n25869), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26022), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_33.INIT1 = 16'h0000;
    defparam count_2613_add_4_33.INJECT1_0 = "NO";
    defparam count_2613_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26021), .COUT(n26022), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_31.INJECT1_0 = "NO";
    defparam count_2613_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25867), .COUT(n25868), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25866), .COUT(n25867), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26020), .COUT(n26021), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_29.INJECT1_0 = "NO";
    defparam count_2613_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26019), .COUT(n26020), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_27.INJECT1_0 = "NO";
    defparam count_2613_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26018), .COUT(n26019), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_25.INJECT1_0 = "NO";
    defparam count_2613_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25865), .COUT(n25866), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25864), .COUT(n25865), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26017), .COUT(n26018), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_23.INJECT1_0 = "NO";
    defparam count_2613_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26016), .COUT(n26017), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_21.INJECT1_0 = "NO";
    defparam count_2613_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25863), .COUT(n25864), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26015), .COUT(n26016), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_19.INJECT1_0 = "NO";
    defparam count_2613_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25862), .COUT(n25863), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26014), .COUT(n26015), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_17.INJECT1_0 = "NO";
    defparam count_2613_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26013), .COUT(n26014), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_15.INJECT1_0 = "NO";
    defparam count_2613_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25861), .COUT(n25862), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25860), .COUT(n25861), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26012), .COUT(n26013), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_13.INJECT1_0 = "NO";
    defparam count_2613_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25859), .COUT(n25860), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26011), .COUT(n26012), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_11.INJECT1_0 = "NO";
    defparam count_2613_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26010), .COUT(n26011), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_9.INJECT1_0 = "NO";
    defparam count_2613_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26009), .COUT(n26010), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_7.INJECT1_0 = "NO";
    defparam count_2613_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25858), .COUT(n25859), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    FD1S3IX count_2613__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i0.GSR = "ENABLED";
    CCU2D count_2613_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26008), .COUT(n26009), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_5.INJECT1_0 = "NO";
    defparam count_2613_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26007), .COUT(n26008), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2613_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2613_add_4_3.INJECT1_0 = "NO";
    defparam count_2613_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2613_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26007), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613_add_4_1.INIT0 = 16'hF000;
    defparam count_2613_add_4_1.INIT1 = 16'h0555;
    defparam count_2613_add_4_1.INJECT1_0 = "NO";
    defparam count_2613_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25857), .COUT(n25858), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25856), .COUT(n25857), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25855), .COUT(n25856), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25855), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25702), .S1(n7851));
    defparam sub_2024_add_2_33.INIT0 = 16'h5555;
    defparam sub_2024_add_2_33.INIT1 = 16'h0000;
    defparam sub_2024_add_2_33.INJECT1_0 = "NO";
    defparam sub_2024_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25701), .COUT(n25702));
    defparam sub_2024_add_2_31.INIT0 = 16'h5999;
    defparam sub_2024_add_2_31.INIT1 = 16'h5999;
    defparam sub_2024_add_2_31.INJECT1_0 = "NO";
    defparam sub_2024_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25700), .COUT(n25701));
    defparam sub_2024_add_2_29.INIT0 = 16'h5999;
    defparam sub_2024_add_2_29.INIT1 = 16'h5999;
    defparam sub_2024_add_2_29.INJECT1_0 = "NO";
    defparam sub_2024_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25699), .COUT(n25700));
    defparam sub_2024_add_2_27.INIT0 = 16'h5999;
    defparam sub_2024_add_2_27.INIT1 = 16'h5999;
    defparam sub_2024_add_2_27.INJECT1_0 = "NO";
    defparam sub_2024_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25698), .COUT(n25699));
    defparam sub_2024_add_2_25.INIT0 = 16'h5999;
    defparam sub_2024_add_2_25.INIT1 = 16'h5999;
    defparam sub_2024_add_2_25.INJECT1_0 = "NO";
    defparam sub_2024_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25697), .COUT(n25698));
    defparam sub_2024_add_2_23.INIT0 = 16'h5999;
    defparam sub_2024_add_2_23.INIT1 = 16'h5999;
    defparam sub_2024_add_2_23.INJECT1_0 = "NO";
    defparam sub_2024_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25696), .COUT(n25697));
    defparam sub_2024_add_2_21.INIT0 = 16'h5999;
    defparam sub_2024_add_2_21.INIT1 = 16'h5999;
    defparam sub_2024_add_2_21.INJECT1_0 = "NO";
    defparam sub_2024_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25695), .COUT(n25696));
    defparam sub_2024_add_2_19.INIT0 = 16'h5999;
    defparam sub_2024_add_2_19.INIT1 = 16'h5999;
    defparam sub_2024_add_2_19.INJECT1_0 = "NO";
    defparam sub_2024_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25694), .COUT(n25695));
    defparam sub_2024_add_2_17.INIT0 = 16'h5999;
    defparam sub_2024_add_2_17.INIT1 = 16'h5999;
    defparam sub_2024_add_2_17.INJECT1_0 = "NO";
    defparam sub_2024_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25693), .COUT(n25694));
    defparam sub_2024_add_2_15.INIT0 = 16'h5999;
    defparam sub_2024_add_2_15.INIT1 = 16'h5999;
    defparam sub_2024_add_2_15.INJECT1_0 = "NO";
    defparam sub_2024_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25692), .COUT(n25693));
    defparam sub_2024_add_2_13.INIT0 = 16'h5999;
    defparam sub_2024_add_2_13.INIT1 = 16'h5999;
    defparam sub_2024_add_2_13.INJECT1_0 = "NO";
    defparam sub_2024_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25691), .COUT(n25692));
    defparam sub_2024_add_2_11.INIT0 = 16'h5999;
    defparam sub_2024_add_2_11.INIT1 = 16'h5999;
    defparam sub_2024_add_2_11.INJECT1_0 = "NO";
    defparam sub_2024_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25690), .COUT(n25691));
    defparam sub_2024_add_2_9.INIT0 = 16'h5999;
    defparam sub_2024_add_2_9.INIT1 = 16'h5999;
    defparam sub_2024_add_2_9.INJECT1_0 = "NO";
    defparam sub_2024_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25689), .COUT(n25690));
    defparam sub_2024_add_2_7.INIT0 = 16'h5999;
    defparam sub_2024_add_2_7.INIT1 = 16'h5999;
    defparam sub_2024_add_2_7.INJECT1_0 = "NO";
    defparam sub_2024_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25688), .COUT(n25689));
    defparam sub_2024_add_2_5.INIT0 = 16'h5999;
    defparam sub_2024_add_2_5.INIT1 = 16'h5999;
    defparam sub_2024_add_2_5.INJECT1_0 = "NO";
    defparam sub_2024_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2024_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25687), .COUT(n25688));
    defparam sub_2024_add_2_3.INIT0 = 16'h5999;
    defparam sub_2024_add_2_3.INIT1 = 16'h5999;
    defparam sub_2024_add_2_3.INJECT1_0 = "NO";
    defparam sub_2024_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n30301), .PD(n16222), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2024_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n25687));
    defparam sub_2024_add_2_1.INIT0 = 16'h0000;
    defparam sub_2024_add_2_1.INIT1 = 16'h5999;
    defparam sub_2024_add_2_1.INJECT1_0 = "NO";
    defparam sub_2024_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25686), .S1(n7886));
    defparam sub_2026_add_2_33.INIT0 = 16'h5999;
    defparam sub_2026_add_2_33.INIT1 = 16'h0000;
    defparam sub_2026_add_2_33.INJECT1_0 = "NO";
    defparam sub_2026_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25685), .COUT(n25686));
    defparam sub_2026_add_2_31.INIT0 = 16'h5999;
    defparam sub_2026_add_2_31.INIT1 = 16'h5999;
    defparam sub_2026_add_2_31.INJECT1_0 = "NO";
    defparam sub_2026_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25684), .COUT(n25685));
    defparam sub_2026_add_2_29.INIT0 = 16'h5999;
    defparam sub_2026_add_2_29.INIT1 = 16'h5999;
    defparam sub_2026_add_2_29.INJECT1_0 = "NO";
    defparam sub_2026_add_2_29.INJECT1_1 = "NO";
    FD1S3IX count_2613__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i1.GSR = "ENABLED";
    CCU2D sub_2026_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25683), .COUT(n25684));
    defparam sub_2026_add_2_27.INIT0 = 16'h5999;
    defparam sub_2026_add_2_27.INIT1 = 16'h5999;
    defparam sub_2026_add_2_27.INJECT1_0 = "NO";
    defparam sub_2026_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25682), .COUT(n25683));
    defparam sub_2026_add_2_25.INIT0 = 16'h5999;
    defparam sub_2026_add_2_25.INIT1 = 16'h5999;
    defparam sub_2026_add_2_25.INJECT1_0 = "NO";
    defparam sub_2026_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25681), .COUT(n25682));
    defparam sub_2026_add_2_23.INIT0 = 16'h5999;
    defparam sub_2026_add_2_23.INIT1 = 16'h5999;
    defparam sub_2026_add_2_23.INJECT1_0 = "NO";
    defparam sub_2026_add_2_23.INJECT1_1 = "NO";
    FD1S3IX count_2613__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i2.GSR = "ENABLED";
    FD1S3IX count_2613__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i3.GSR = "ENABLED";
    FD1S3IX count_2613__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i4.GSR = "ENABLED";
    FD1S3IX count_2613__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i5.GSR = "ENABLED";
    FD1S3IX count_2613__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i6.GSR = "ENABLED";
    FD1S3IX count_2613__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i7.GSR = "ENABLED";
    FD1S3IX count_2613__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i8.GSR = "ENABLED";
    FD1S3IX count_2613__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i9.GSR = "ENABLED";
    FD1S3IX count_2613__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i10.GSR = "ENABLED";
    FD1S3IX count_2613__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i11.GSR = "ENABLED";
    FD1S3IX count_2613__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i12.GSR = "ENABLED";
    FD1S3IX count_2613__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i13.GSR = "ENABLED";
    FD1S3IX count_2613__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i14.GSR = "ENABLED";
    FD1S3IX count_2613__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i15.GSR = "ENABLED";
    FD1S3IX count_2613__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i16.GSR = "ENABLED";
    FD1S3IX count_2613__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i17.GSR = "ENABLED";
    FD1S3IX count_2613__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i18.GSR = "ENABLED";
    FD1S3IX count_2613__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i19.GSR = "ENABLED";
    FD1S3IX count_2613__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i20.GSR = "ENABLED";
    FD1S3IX count_2613__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i21.GSR = "ENABLED";
    FD1S3IX count_2613__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i22.GSR = "ENABLED";
    FD1S3IX count_2613__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i23.GSR = "ENABLED";
    FD1S3IX count_2613__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i24.GSR = "ENABLED";
    FD1S3IX count_2613__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i25.GSR = "ENABLED";
    FD1S3IX count_2613__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i26.GSR = "ENABLED";
    FD1S3IX count_2613__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i27.GSR = "ENABLED";
    FD1S3IX count_2613__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i28.GSR = "ENABLED";
    FD1S3IX count_2613__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i29.GSR = "ENABLED";
    FD1S3IX count_2613__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i30.GSR = "ENABLED";
    FD1S3IX count_2613__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n30301), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2613__i31.GSR = "ENABLED";
    CCU2D sub_2026_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25680), .COUT(n25681));
    defparam sub_2026_add_2_21.INIT0 = 16'h5999;
    defparam sub_2026_add_2_21.INIT1 = 16'h5999;
    defparam sub_2026_add_2_21.INJECT1_0 = "NO";
    defparam sub_2026_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25679), .COUT(n25680));
    defparam sub_2026_add_2_19.INIT0 = 16'h5999;
    defparam sub_2026_add_2_19.INIT1 = 16'h5999;
    defparam sub_2026_add_2_19.INJECT1_0 = "NO";
    defparam sub_2026_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25678), .COUT(n25679));
    defparam sub_2026_add_2_17.INIT0 = 16'h5999;
    defparam sub_2026_add_2_17.INIT1 = 16'h5999;
    defparam sub_2026_add_2_17.INJECT1_0 = "NO";
    defparam sub_2026_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25677), .COUT(n25678));
    defparam sub_2026_add_2_15.INIT0 = 16'h5999;
    defparam sub_2026_add_2_15.INIT1 = 16'h5999;
    defparam sub_2026_add_2_15.INJECT1_0 = "NO";
    defparam sub_2026_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25676), .COUT(n25677));
    defparam sub_2026_add_2_13.INIT0 = 16'h5999;
    defparam sub_2026_add_2_13.INIT1 = 16'h5999;
    defparam sub_2026_add_2_13.INJECT1_0 = "NO";
    defparam sub_2026_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25675), .COUT(n25676));
    defparam sub_2026_add_2_11.INIT0 = 16'h5999;
    defparam sub_2026_add_2_11.INIT1 = 16'h5999;
    defparam sub_2026_add_2_11.INJECT1_0 = "NO";
    defparam sub_2026_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25674), .COUT(n25675));
    defparam sub_2026_add_2_9.INIT0 = 16'h5999;
    defparam sub_2026_add_2_9.INIT1 = 16'h5999;
    defparam sub_2026_add_2_9.INJECT1_0 = "NO";
    defparam sub_2026_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25673), .COUT(n25674));
    defparam sub_2026_add_2_7.INIT0 = 16'h5999;
    defparam sub_2026_add_2_7.INIT1 = 16'h5999;
    defparam sub_2026_add_2_7.INJECT1_0 = "NO";
    defparam sub_2026_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n30301), .CD(n16222), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2026_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25672), .COUT(n25673));
    defparam sub_2026_add_2_5.INIT0 = 16'h5999;
    defparam sub_2026_add_2_5.INIT1 = 16'h5999;
    defparam sub_2026_add_2_5.INJECT1_0 = "NO";
    defparam sub_2026_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25671), .COUT(n25672));
    defparam sub_2026_add_2_3.INIT0 = 16'h5999;
    defparam sub_2026_add_2_3.INIT1 = 16'h5999;
    defparam sub_2026_add_2_3.INJECT1_0 = "NO";
    defparam sub_2026_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2026_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n25671));
    defparam sub_2026_add_2_1.INIT0 = 16'h0000;
    defparam sub_2026_add_2_1.INIT1 = 16'h5999;
    defparam sub_2026_add_2_1.INJECT1_0 = "NO";
    defparam sub_2026_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25670), .S1(n7920));
    defparam sub_2027_add_2_33.INIT0 = 16'hf555;
    defparam sub_2027_add_2_33.INIT1 = 16'h0000;
    defparam sub_2027_add_2_33.INJECT1_0 = "NO";
    defparam sub_2027_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25669), .COUT(n25670));
    defparam sub_2027_add_2_31.INIT0 = 16'hf555;
    defparam sub_2027_add_2_31.INIT1 = 16'hf555;
    defparam sub_2027_add_2_31.INJECT1_0 = "NO";
    defparam sub_2027_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25668), .COUT(n25669));
    defparam sub_2027_add_2_29.INIT0 = 16'hf555;
    defparam sub_2027_add_2_29.INIT1 = 16'hf555;
    defparam sub_2027_add_2_29.INJECT1_0 = "NO";
    defparam sub_2027_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25667), .COUT(n25668));
    defparam sub_2027_add_2_27.INIT0 = 16'hf555;
    defparam sub_2027_add_2_27.INIT1 = 16'hf555;
    defparam sub_2027_add_2_27.INJECT1_0 = "NO";
    defparam sub_2027_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25666), .COUT(n25667));
    defparam sub_2027_add_2_25.INIT0 = 16'hf555;
    defparam sub_2027_add_2_25.INIT1 = 16'hf555;
    defparam sub_2027_add_2_25.INJECT1_0 = "NO";
    defparam sub_2027_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25665), .COUT(n25666));
    defparam sub_2027_add_2_23.INIT0 = 16'hf555;
    defparam sub_2027_add_2_23.INIT1 = 16'hf555;
    defparam sub_2027_add_2_23.INJECT1_0 = "NO";
    defparam sub_2027_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25664), .COUT(n25665));
    defparam sub_2027_add_2_21.INIT0 = 16'hf555;
    defparam sub_2027_add_2_21.INIT1 = 16'hf555;
    defparam sub_2027_add_2_21.INJECT1_0 = "NO";
    defparam sub_2027_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25663), .COUT(n25664));
    defparam sub_2027_add_2_19.INIT0 = 16'hf555;
    defparam sub_2027_add_2_19.INIT1 = 16'hf555;
    defparam sub_2027_add_2_19.INJECT1_0 = "NO";
    defparam sub_2027_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25662), .COUT(n25663));
    defparam sub_2027_add_2_17.INIT0 = 16'hf555;
    defparam sub_2027_add_2_17.INIT1 = 16'hf555;
    defparam sub_2027_add_2_17.INJECT1_0 = "NO";
    defparam sub_2027_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25661), .COUT(n25662));
    defparam sub_2027_add_2_15.INIT0 = 16'hf555;
    defparam sub_2027_add_2_15.INIT1 = 16'hf555;
    defparam sub_2027_add_2_15.INJECT1_0 = "NO";
    defparam sub_2027_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2027_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25660), .COUT(n25661));
    defparam sub_2027_add_2_13.INIT0 = 16'hf555;
    defparam sub_2027_add_2_13.INIT1 = 16'hf555;
    defparam sub_2027_add_2_13.INJECT1_0 = "NO";
    defparam sub_2027_add_2_13.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module SabertoothSerialPeripheral
//

module SabertoothSerialPeripheral (debug_c_c, n9122, n282, n32384, \databus[6] , 
            \databus[5] , \databus[4] , \databus[3] , \databus[2] , 
            \databus[1] , \databus[0] , n32385, \read_size[0] , n21563, 
            n32381, \select[2] , \register_addr[0] , n30422, \register_addr[1] , 
            \register_addr[3] , \register_addr[2] , n30445, n32380, 
            rw, n5, n5_adj_221, n5_adj_222, n5_adj_223, n5_adj_224, 
            n5_adj_225, n5_adj_226, n5_adj_227, n30488, n13269, n30350, 
            n30314, n30324, n13534, n30349, n30491, n30489, n30379, 
            n28137, n30478, n8, \state[0] , GND_net, n12, n30305, 
            n31, n27462, n22, n19, n32382, \reset_count[14] , \reset_count[12] , 
            n28605, motor_pwm_l_c, n30342, select_clk, n107, n8129) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n9122;
    input n282;
    input n32384;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    input \databus[0] ;
    input n32385;
    output \read_size[0] ;
    output n21563;
    input n32381;
    input \select[2] ;
    input \register_addr[0] ;
    input n30422;
    input \register_addr[1] ;
    input \register_addr[3] ;
    input \register_addr[2] ;
    output n30445;
    input n32380;
    input rw;
    output n5;
    output n5_adj_221;
    output n5_adj_222;
    output n5_adj_223;
    output n5_adj_224;
    output n5_adj_225;
    output n5_adj_226;
    output n5_adj_227;
    input n30488;
    input n13269;
    input n30350;
    output n30314;
    input n30324;
    output n13534;
    input n30349;
    input n30491;
    input n30489;
    output n30379;
    output n28137;
    input n30478;
    output n8;
    output \state[0] ;
    input GND_net;
    input n12;
    input n30305;
    output n31;
    input n27462;
    output n22;
    input n19;
    input n32382;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input n28605;
    output motor_pwm_l_c;
    input n30342;
    output select_clk;
    input n107;
    output n8129;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [7:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(92[12:22])
    
    wire n2635;
    wire [7:0]n28;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n13546, n30323;
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n21773, n30322, prev_select;
    wire [7:0]n27;
    
    wire n30526, n30525, n26372, n9032, n28510;
    
    FD1P3IX read_value__i7 (.D(n28[7]), .SP(n2635), .CD(n9122), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n28[6]), .SP(n2635), .CD(n9122), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n28[5]), .SP(n2635), .CD(n9122), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n28[4]), .SP(n2635), .CD(n9122), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n28[3]), .SP(n2635), .CD(n9122), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX register_0__i16 (.D(n282), .SP(n13546), .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n30323), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n30323), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n30323), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n30323), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n30323), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n30323), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n30323), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n282), .SP(n21773), .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n30322), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n30322), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n30322), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n30322), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n30322), .PD(n32384), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n30322), .PD(n32385), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i2.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n28[2]), .SP(n2635), .CD(n9122), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n21563), .SP(n2635), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n30322), .PD(n32381), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam prev_select_138.GSR = "ENABLED";
    LUT4 mux_1881_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n28[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1881_Mux_7_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n28[0]), .SP(n2635), .CD(n9122), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3AX read_value__i1 (.D(n27[1]), .SP(n2635), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1881_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n28[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1881_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1881_Mux_2_i1_3_lut (.A(\register[0] [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n28[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1881_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1881_Mux_5_i1_3_lut (.A(\register[0] [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n28[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1881_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_3_lut_4_lut_then_4_lut (.A(n30422), .B(\register_addr[1] ), 
         .C(\register_addr[3] ), .D(\register_addr[2] ), .Z(n30526)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_3_lut_3_lut_4_lut_then_4_lut.init = 16'h0004;
    LUT4 i1_3_lut_3_lut_4_lut_else_4_lut (.A(n30422), .B(\register_addr[3] ), 
         .C(\register_addr[2] ), .Z(n30525)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i1_3_lut_3_lut_4_lut_else_4_lut.init = 16'h0101;
    LUT4 i1_2_lut_rep_436 (.A(\select[2] ), .B(prev_select), .Z(n30445)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_rep_436.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\select[2] ), .B(prev_select), .C(n32380), 
         .Z(n2635)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 mux_1881_Mux_4_i1_3_lut (.A(\register[0] [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n28[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1881_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 Select_4227_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[0]), 
         .Z(n5)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4227_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4226_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[1]), 
         .Z(n5_adj_221)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4226_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4224_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[3]), 
         .Z(n5_adj_222)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4224_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4225_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[2]), 
         .Z(n5_adj_223)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4225_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4223_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[4]), 
         .Z(n5_adj_224)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4223_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4222_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[5]), 
         .Z(n5_adj_225)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4222_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4221_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[6]), 
         .Z(n5_adj_226)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4221_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4220_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[7]), 
         .Z(n5_adj_227)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4220_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 i21695_3_lut_rep_305_4_lut_4_lut (.A(n30488), .B(n13269), .C(n30350), 
         .D(rw), .Z(n30314)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i21695_3_lut_rep_305_4_lut_4_lut.init = 16'h0010;
    LUT4 i21729_2_lut_4_lut_4_lut (.A(n30488), .B(n32380), .C(n13269), 
         .D(n30324), .Z(n13534)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i21729_2_lut_4_lut_4_lut.init = 16'hcdcc;
    LUT4 mux_1881_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n28[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1881_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1881_Mux_3_i1_3_lut (.A(\register[0] [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n28[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1881_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 i14960_4_lut (.A(\register[0] [1]), .B(n9122), .C(\register[1] [1]), 
         .D(\register_addr[0] ), .Z(n27[1])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam i14960_4_lut.init = 16'h3022;
    LUT4 i21732_2_lut_3_lut (.A(\register_addr[0] ), .B(n30349), .C(n32380), 
         .Z(n21773)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(131[9] 136[16])
    defparam i21732_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i2_2_lut_rep_370_3_lut_4_lut (.A(n30491), .B(n30488), .C(n30489), 
         .D(\register_addr[1] ), .Z(n30379)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i2_2_lut_rep_370_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21670_2_lut_2_lut_3_lut_4_lut (.A(n30491), .B(n30488), .C(\register_addr[1] ), 
         .D(n30489), .Z(n21563)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i21670_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n30491), .B(n30488), .C(\register_addr[1] ), 
         .D(n30489), .Z(n28137)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n30349), .C(n32380), 
         .Z(n13546)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(131[9] 136[16])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut_4_lut (.A(\register[0] [7]), .B(n30478), .C(\register[0] [1]), 
         .D(n26372), .Z(n9032)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h2000;
    LUT4 i21362_3_lut_4_lut_4_lut (.A(\register[0] [7]), .B(n30478), .C(\register[0] [1]), 
         .D(n26372), .Z(n28510)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i21362_3_lut_4_lut_4_lut.init = 16'heccc;
    LUT4 i21691_2_lut_rep_313_4_lut (.A(rw), .B(n30445), .C(n30379), .D(\register_addr[0] ), 
         .Z(n30322)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i21691_2_lut_rep_313_4_lut.init = 16'h0004;
    LUT4 i4499_2_lut_rep_314_4_lut (.A(rw), .B(n30445), .C(n30379), .D(\register_addr[0] ), 
         .Z(n30323)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i4499_2_lut_rep_314_4_lut.init = 16'h0400;
    PFUMX i22351 (.BLUT(n30525), .ALUT(n30526), .C0(\register_addr[0] ), 
          .Z(n8));
    SabertoothSerial sserial (.\register[0][3] (\register[0] [3]), .n9032(n9032), 
            .n30478(n30478), .\register[1][3] (\register[1] [3]), .\register[1][7] (\register[1] [7]), 
            .\register[1][1] (\register[1] [1]), .\register[0][4] (\register[0] [4]), 
            .\register[0][2] (\register[0] [2]), .n26372(n26372), .\register[0][5] (\register[0] [5]), 
            .\register[0][6] (\register[0] [6]), .\register[1][4] (\register[1] [4]), 
            .\register[1][5] (\register[1] [5]), .\register[1][2] (\register[1] [2]), 
            .\state[0] (\state[0] ), .debug_c_c(debug_c_c), .GND_net(GND_net), 
            .n12(n12), .n30305(n30305), .n31(n31), .n27462(n27462), 
            .n22(n22), .\register[1][6] (\register[1] [6]), .\register[0][1] (\register[0] [1]), 
            .\register[0][7] (\register[0] [7]), .n28510(n28510), .n19(n19), 
            .n32382(n32382), .\reset_count[14] (\reset_count[14] ), .\reset_count[12] (\reset_count[12] ), 
            .n28605(n28605), .n32380(n32380), .motor_pwm_l_c(motor_pwm_l_c), 
            .n30342(n30342), .select_clk(select_clk), .n107(n107), .n8129(n8129)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(142[19] 147[34])
    
endmodule
//
// Verilog Description of module SabertoothSerial
//

module SabertoothSerial (\register[0][3] , n9032, n30478, \register[1][3] , 
            \register[1][7] , \register[1][1] , \register[0][4] , \register[0][2] , 
            n26372, \register[0][5] , \register[0][6] , \register[1][4] , 
            \register[1][5] , \register[1][2] , \state[0] , debug_c_c, 
            GND_net, n12, n30305, n31, n27462, n22, \register[1][6] , 
            \register[0][1] , \register[0][7] , n28510, n19, n32382, 
            \reset_count[14] , \reset_count[12] , n28605, n32380, motor_pwm_l_c, 
            n30342, select_clk, n107, n8129) /* synthesis syn_module_defined=1 */ ;
    input \register[0][3] ;
    input n9032;
    input n30478;
    input \register[1][3] ;
    input \register[1][7] ;
    input \register[1][1] ;
    input \register[0][4] ;
    input \register[0][2] ;
    output n26372;
    input \register[0][5] ;
    input \register[0][6] ;
    input \register[1][4] ;
    input \register[1][5] ;
    input \register[1][2] ;
    output \state[0] ;
    input debug_c_c;
    input GND_net;
    input n12;
    input n30305;
    output n31;
    input n27462;
    output n22;
    input \register[1][6] ;
    input \register[0][1] ;
    input \register[0][7] ;
    input n28510;
    input n19;
    input n32382;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input n28605;
    input n32380;
    output motor_pwm_l_c;
    input n30342;
    output select_clk;
    input n107;
    output n8129;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30476;
    wire [31:0]n17;
    
    wire n9035, n30477;
    wire [31:0]n63;
    
    wire n30423, n6, n28176;
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    wire [3:0]n16;
    
    wire n17845, n29, n26, n24, n29_adj_492, n26_adj_493, n24_adj_494, 
        n29_adj_495, n26_adj_496, n36, n30, n28, n21, n27999, 
        n30_adj_497, n36_adj_498, n30_adj_499, n28_adj_500;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(16[12:19])
    
    wire n30304, n27, n24_adj_501, n977, n30460, n30419, n30341, 
        n27456;
    wire [7:0]n5312;
    
    wire n27360, n27302, n27116, n27300, n30418, n30390, n30389, 
        n12238, n30365, n7;
    
    LUT4 i15041_4_lut (.A(\register[0][3] ), .B(n9032), .C(n30478), .D(n30476), 
         .Z(n17[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(37[20:73])
    defparam i15041_4_lut.init = 16'hcdce;
    LUT4 i15046_4_lut (.A(\register[1][3] ), .B(n9035), .C(n30478), .D(n30477), 
         .Z(n63[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15046_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut (.A(\register[1][7] ), .B(n30478), .C(n30423), .D(\register[1][1] ), 
         .Z(n9035)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h2000;
    LUT4 i4_4_lut (.A(\register[0][4] ), .B(\register[0][2] ), .C(\register[0][3] ), 
         .D(n6), .Z(n26372)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(\register[0][5] ), .B(\register[0][6] ), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i3_4_lut (.A(\register[1][4] ), .B(\register[1][3] ), .C(\register[1][5] ), 
         .D(\register[1][2] ), .Z(n28176)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    FD1S3IX state__i0 (.D(n12), .CK(debug_c_c), .CD(GND_net), .Q(\state[0] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3IX state__i1 (.D(n16[1]), .SP(n30305), .CD(GND_net), .CK(debug_c_c), 
            .Q(state[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i1.GSR = "ENABLED";
    PFUMX i11436 (.BLUT(n17[2]), .ALUT(n63[2]), .C0(state[1]), .Z(n17845));
    PFUMX i39 (.BLUT(n29), .ALUT(n26), .C0(state[1]), .Z(n24));
    PFUMX i39_adj_383 (.BLUT(n29_adj_492), .ALUT(n26_adj_493), .C0(state[1]), 
          .Z(n24_adj_494));
    PFUMX i44 (.BLUT(n29_adj_495), .ALUT(n26_adj_496), .C0(state[1]), 
          .Z(n31));
    PFUMX i48 (.BLUT(n36), .ALUT(n30), .C0(state[1]), .Z(n28));
    PFUMX i38 (.BLUT(n21), .ALUT(n27999), .C0(state[1]), .Z(n30_adj_497));
    PFUMX i48_adj_384 (.BLUT(n36_adj_498), .ALUT(n30_adj_499), .C0(state[1]), 
          .Z(n28_adj_500));
    FD1P3AX tx_data_i0_i0 (.D(n27462), .SP(n30304), .CK(debug_c_c), .Q(tx_data[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    PFUMX i35 (.BLUT(n27), .ALUT(n24_adj_501), .C0(state[1]), .Z(n22));
    FD1P3AX send_31 (.D(n30460), .SP(n30305), .CK(debug_c_c), .Q(n977));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam send_31.GSR = "ENABLED";
    LUT4 i21331_2_lut_rep_332_3_lut_4_lut (.A(\register[1][4] ), .B(n30419), 
         .C(\register[1][6] ), .D(\register[1][5] ), .Z(n30341)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i21331_2_lut_rep_332_3_lut_4_lut.init = 16'h8000;
    LUT4 i6_1_lut_rep_451 (.A(\state[0] ), .Z(n30460)) /* synthesis lut_function=(!(A)) */ ;
    defparam i6_1_lut_rep_451.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(\state[0] ), .B(n24), .Z(n27456)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_385 (.A(\state[0] ), .B(n17845), .Z(n5312[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_385.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_386 (.A(\state[0] ), .B(n24_adj_494), .Z(n27360)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_386.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_387 (.A(\state[0] ), .B(n28_adj_500), .Z(n27302)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_387.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_388 (.A(\state[0] ), .B(n28), .Z(n27116)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_388.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_389 (.A(\state[0] ), .B(n30_adj_497), .Z(n27300)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_389.init = 16'h4444;
    LUT4 i1_4_lut_adj_390 (.A(n9032), .B(n30478), .C(\register[0][1] ), 
         .D(\register[0][2] ), .Z(n29)) /* synthesis lut_function=(A+!(B+(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_390.init = 16'habba;
    LUT4 i1_4_lut_adj_391 (.A(n30478), .B(n9035), .C(\register[1][2] ), 
         .D(\register[1][1] ), .Z(n26)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_391.init = 16'hcddc;
    LUT4 i9_2_lut (.A(state[1]), .B(\state[0] ), .Z(n16[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    defparam i9_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_392 (.A(n9032), .B(n30478), .C(n30418), .D(\register[0][4] ), 
         .Z(n29_adj_492)) /* synthesis lut_function=(A+!(B+(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_392.init = 16'habba;
    LUT4 i1_4_lut_adj_393 (.A(n30478), .B(n9035), .C(\register[1][4] ), 
         .D(n30419), .Z(n26_adj_493)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_393.init = 16'hcddc;
    LUT4 i5139_2_lut_rep_467 (.A(\register[0][2] ), .B(\register[0][1] ), 
         .Z(n30476)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5139_2_lut_rep_467.init = 16'h8888;
    LUT4 i5825_2_lut_rep_381_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n30390)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5825_2_lut_rep_381_3_lut_4_lut.init = 16'h8000;
    LUT4 i5141_2_lut_rep_409_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n30418)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5141_2_lut_rep_409_3_lut.init = 16'h8080;
    LUT4 i4735_2_lut_rep_468 (.A(\register[1][2] ), .B(\register[1][1] ), 
         .Z(n30477)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4735_2_lut_rep_468.init = 16'h8888;
    LUT4 i5785_2_lut_rep_380_3_lut_4_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][4] ), .D(\register[1][3] ), .Z(n30389)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5785_2_lut_rep_380_3_lut_4_lut.init = 16'h8000;
    LUT4 i4828_2_lut_rep_410_3_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][3] ), .Z(n30419)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i4828_2_lut_rep_410_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_394 (.A(n9032), .B(\register[0][7] ), .C(\register[0][6] ), 
         .D(n12238), .Z(n29_adj_495)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C (D))))) */ ;
    defparam i1_4_lut_adj_394.init = 16'h4111;
    LUT4 i1_3_lut_4_lut (.A(n30365), .B(\register[1][6] ), .C(\register[1][7] ), 
         .D(n9035), .Z(n26_adj_496)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A (C+(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0087;
    LUT4 i5827_2_lut_3_lut_4_lut (.A(\register[0][3] ), .B(n30476), .C(\register[0][5] ), 
         .D(\register[0][4] ), .Z(n12238)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5827_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i5819_2_lut_rep_356_3_lut_4_lut (.A(\register[1][3] ), .B(n30477), 
         .C(\register[1][5] ), .D(\register[1][4] ), .Z(n30365)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5819_2_lut_rep_356_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_414 (.A(\register[1][6] ), .B(n28176), .Z(n30423)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_414.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_395 (.A(\register[1][6] ), .B(n28176), .C(\register[1][7] ), 
         .D(\register[1][1] ), .Z(n24_adj_501)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i1_3_lut_4_lut_adj_395.init = 16'h80ff;
    LUT4 i1_4_lut_adj_396 (.A(n9032), .B(n30478), .C(n12238), .D(\register[0][6] ), 
         .Z(n36)) /* synthesis lut_function=(A+!(B+(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_396.init = 16'habba;
    LUT4 i1_4_lut_adj_397 (.A(n9035), .B(n30478), .C(n30365), .D(\register[1][6] ), 
         .Z(n30)) /* synthesis lut_function=(A+!(B+(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_397.init = 16'habba;
    LUT4 i4_4_lut_adj_398 (.A(n28510), .B(n12238), .C(\register[0][6] ), 
         .D(\register[0][7] ), .Z(n21)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i4_4_lut_adj_398.init = 16'h4000;
    LUT4 i1_4_lut_adj_399 (.A(n30478), .B(\register[1][7] ), .C(n30341), 
         .D(n7), .Z(n27999)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_399.init = 16'hffbf;
    LUT4 i1_2_lut_adj_400 (.A(\register[1][1] ), .B(n28176), .Z(n7)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_400.init = 16'h8888;
    FD1P3AX tx_data_i0_i1 (.D(n27456), .SP(n30304), .CK(debug_c_c), .Q(tx_data[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i2 (.D(n5312[2]), .SP(n30304), .CK(debug_c_c), 
            .Q(tx_data[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n27360), .SP(n30304), .CK(debug_c_c), .Q(tx_data[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n27302), .SP(n30304), .CK(debug_c_c), .Q(tx_data[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i5 (.D(n27116), .SP(n30304), .CK(debug_c_c), .Q(tx_data[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i6 (.D(n19), .SP(n30304), .CK(debug_c_c), .Q(tx_data[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i7 (.D(n27300), .SP(n30304), .CK(debug_c_c), .Q(tx_data[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_401 (.A(n9032), .B(n30478), .C(n30390), .D(\register[0][5] ), 
         .Z(n36_adj_498)) /* synthesis lut_function=(A+!(B+(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_401.init = 16'habba;
    LUT4 i1_4_lut_adj_402 (.A(n9035), .B(n30478), .C(n30389), .D(\register[1][5] ), 
         .Z(n30_adj_499)) /* synthesis lut_function=(A+!(B+(C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_402.init = 16'habba;
    LUT4 i1_3_lut (.A(\register[0][7] ), .B(\register[0][1] ), .C(n26372), 
         .Z(n27)) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;
    defparam i1_3_lut.init = 16'hb3b3;
    \UARTTransmitter(baud_div=1250)  sender (.n32382(n32382), .n977(n977), 
            .\reset_count[14] (\reset_count[14] ), .\reset_count[12] (\reset_count[12] ), 
            .n28605(n28605), .n32380(n32380), .tx_data({tx_data}), .motor_pwm_l_c(motor_pwm_l_c), 
            .n30342(n30342), .debug_c_c(debug_c_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(63[26] 67[47])
    \ClockDividerP(factor=12000)  baud_gen (.debug_c_c(debug_c_c), .select_clk(select_clk), 
            .n107(n107), .GND_net(GND_net), .n8129(n8129), .\state[0] (\state[0] ), 
            .n32380(n32380), .n30304(n30304)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(21[25] 23[48])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=1250) 
//

module \UARTTransmitter(baud_div=1250)  (n32382, n977, \reset_count[14] , 
            \reset_count[12] , n28605, n32380, tx_data, motor_pwm_l_c, 
            n30342, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    input n32382;
    input n977;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input n28605;
    input n32380;
    input [7:0]tx_data;
    output motor_pwm_l_c;
    input n30342;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n30201, n29690, n7, n10, n104, n30199, n30200, n28054, 
        n9039, n21159, n30315, n2596, n28246, n29651, n14316, 
        n27346, n28634, n28635, n28636;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n28247, n2;
    
    FD1S3IX state__i0 (.D(n30201), .CK(bclk), .CD(n32382), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 state_0__bdd_4_lut (.A(state[0]), .B(state[1]), .C(state[3]), 
         .D(state[2]), .Z(n29690)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam state_0__bdd_4_lut.init = 16'h0f7e;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;
    LUT4 state_2__bdd_2_lut (.A(state[0]), .B(state[3]), .Z(n30199)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_2__bdd_2_lut.init = 16'h1111;
    LUT4 state_2__bdd_4_lut (.A(state[0]), .B(state[3]), .C(n977), .D(state[1]), 
         .Z(n30200)) /* synthesis lut_function=(A (B (C (D)))+!A (B+(C+(D)))) */ ;
    defparam state_2__bdd_4_lut.init = 16'hd554;
    LUT4 i3_4_lut (.A(n977), .B(\reset_count[14] ), .C(state[2]), .D(n28054), 
         .Z(n9039)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i3_4_lut.init = 16'h0800;
    LUT4 i2_4_lut (.A(state[1]), .B(n21159), .C(\reset_count[12] ), .D(n28605), 
         .Z(n28054)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i2_4_lut.init = 16'h1110;
    LUT4 i1_3_lut_rep_306 (.A(n32380), .B(state[2]), .C(state[3]), .Z(n30315)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam i1_3_lut_rep_306.init = 16'h1515;
    LUT4 i1_3_lut_4_lut (.A(n32380), .B(state[2]), .C(state[3]), .D(n2596), 
         .Z(n28246)) /* synthesis lut_function=(!(A+(B (C+(D))+!B !(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1104;
    LUT4 i21811_3_lut (.A(n32380), .B(n29651), .C(state[2]), .Z(n14316)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i21811_3_lut.init = 16'hfbfb;
    LUT4 n977_bdd_4_lut (.A(n977), .B(state[1]), .C(state[3]), .D(state[0]), 
         .Z(n29651)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam n977_bdd_4_lut.init = 16'h8001;
    LUT4 i1_4_lut (.A(n32380), .B(state[3]), .C(state[2]), .D(n2596), 
         .Z(n27346)) /* synthesis lut_function=(!(A+(B (C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h1404;
    LUT4 i916_2_lut (.A(state[0]), .B(state[1]), .Z(n2596)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i916_2_lut.init = 16'h8888;
    PFUMX i21483 (.BLUT(n28634), .ALUT(n28635), .C0(state[1]), .Z(n28636));
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9039), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    FD1P3AX state__i3 (.D(n27346), .SP(n14316), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(state[1]), .B(n30315), .C(state[0]), .Z(n28247)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    PFUMX i22270 (.BLUT(n30200), .ALUT(n30199), .C0(state[2]), .Z(n30201));
    LUT4 i21481_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n28634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21481_3_lut.init = 16'hcaca;
    LUT4 i21482_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n28635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21482_3_lut.init = 16'hcaca;
    LUT4 i14784_2_lut (.A(state[3]), .B(state[0]), .Z(n21159)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14784_2_lut.init = 16'heeee;
    FD1P3AX state__i2 (.D(n28246), .SP(n14316), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n28247), .SP(n14316), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n28636), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    FD1P3JX tx_35 (.D(n104), .SP(n29690), .PD(n30342), .CK(bclk), .Q(motor_pwm_l_c)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15121_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15121_4_lut.init = 16'hfcee;
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9039), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9039), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9039), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9039), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9039), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9039), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9039), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    \ClockDividerP(factor=1250)  baud_gen (.debug_c_c(debug_c_c), .GND_net(GND_net), 
            .bclk(bclk)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=1250) 
//

module \ClockDividerP(factor=1250)  (debug_c_c, GND_net, bclk) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input GND_net;
    output bclk;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n16173;
    wire [31:0]n102;
    
    wire n26150, n26149, n26148, n26147, n26146, n26145, n26144, 
        n26143, n26142, n8164, n26141, n26835, n8, n26140, n39, 
        n52, n48, n40, n31, n50, n44, n32, n26139, n42, n46, 
        n36, n26138, n26137, n26136, n26135, n26261, n26260, n26259, 
        n26258, n26257, n26256, n26255, n26254, n26253, n26252, 
        n26251, n26250, n26249, n26248, n26247;
    
    FD1S3IX count_2618__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i0.GSR = "ENABLED";
    CCU2D count_2618_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26150), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_33.INIT1 = 16'h0000;
    defparam count_2618_add_4_33.INJECT1_0 = "NO";
    defparam count_2618_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26149), .COUT(n26150), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_31.INJECT1_0 = "NO";
    defparam count_2618_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26148), .COUT(n26149), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_29.INJECT1_0 = "NO";
    defparam count_2618_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26147), .COUT(n26148), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_27.INJECT1_0 = "NO";
    defparam count_2618_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26146), .COUT(n26147), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_25.INJECT1_0 = "NO";
    defparam count_2618_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26145), .COUT(n26146), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_23.INJECT1_0 = "NO";
    defparam count_2618_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26144), .COUT(n26145), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_21.INJECT1_0 = "NO";
    defparam count_2618_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26143), .COUT(n26144), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_19.INJECT1_0 = "NO";
    defparam count_2618_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26142), .COUT(n26143), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_17.INJECT1_0 = "NO";
    defparam count_2618_add_4_17.INJECT1_1 = "NO";
    FD1S3AX clk_o_14 (.D(n8164), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2618_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26141), .COUT(n26142), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_15.INJECT1_0 = "NO";
    defparam count_2618_add_4_15.INJECT1_1 = "NO";
    LUT4 i21741_4_lut (.A(n26835), .B(count[5]), .C(n8), .D(count[0]), 
         .Z(n16173)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21741_4_lut.init = 16'h4000;
    CCU2D count_2618_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26140), .COUT(n26141), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_13.INJECT1_0 = "NO";
    defparam count_2618_add_4_13.INJECT1_1 = "NO";
    LUT4 i26_4_lut (.A(n39), .B(n52), .C(n48), .D(n40), .Z(n26835)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i3_3_lut (.A(count[10]), .B(count[6]), .C(count[7]), .Z(n8)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3_3_lut.init = 16'h8080;
    LUT4 i12_2_lut (.A(count[30]), .B(count[13]), .Z(n39)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i12_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(n31), .B(n50), .C(n44), .D(n32), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    CCU2D count_2618_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26139), .COUT(n26140), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_11.INJECT1_0 = "NO";
    defparam count_2618_add_4_11.INJECT1_1 = "NO";
    LUT4 i21_4_lut (.A(count[27]), .B(n42), .C(count[23]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(count[22]), .B(count[18]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i4_2_lut (.A(count[28]), .B(count[9]), .Z(n31)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(count[19]), .B(n46), .C(n36), .D(count[25]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(count[4]), .B(count[11]), .C(count[8]), .D(count[14]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[12]), .B(count[1]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[20]), .B(count[2]), .C(count[24]), .D(count[29]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(count[26]), .B(count[3]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i15_4_lut (.A(count[16]), .B(count[15]), .C(count[31]), .D(count[21]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_4_lut.init = 16'hfffe;
    CCU2D count_2618_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26138), .COUT(n26139), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_9.INJECT1_0 = "NO";
    defparam count_2618_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26137), .COUT(n26138), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_7.INJECT1_0 = "NO";
    defparam count_2618_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26136), .COUT(n26137), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_5.INJECT1_0 = "NO";
    defparam count_2618_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26135), .COUT(n26136), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2618_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2618_add_4_3.INJECT1_0 = "NO";
    defparam count_2618_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2618_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26135), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618_add_4_1.INIT0 = 16'hF000;
    defparam count_2618_add_4_1.INIT1 = 16'h0555;
    defparam count_2618_add_4_1.INJECT1_0 = "NO";
    defparam count_2618_add_4_1.INJECT1_1 = "NO";
    CCU2D add_19123_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26261), 
          .S1(n8164));
    defparam add_19123_32.INIT0 = 16'h5555;
    defparam add_19123_32.INIT1 = 16'h0000;
    defparam add_19123_32.INJECT1_0 = "NO";
    defparam add_19123_32.INJECT1_1 = "NO";
    CCU2D add_19123_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26260), .COUT(n26261));
    defparam add_19123_30.INIT0 = 16'h5555;
    defparam add_19123_30.INIT1 = 16'h5555;
    defparam add_19123_30.INJECT1_0 = "NO";
    defparam add_19123_30.INJECT1_1 = "NO";
    CCU2D add_19123_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26259), .COUT(n26260));
    defparam add_19123_28.INIT0 = 16'h5555;
    defparam add_19123_28.INIT1 = 16'h5555;
    defparam add_19123_28.INJECT1_0 = "NO";
    defparam add_19123_28.INJECT1_1 = "NO";
    CCU2D add_19123_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26258), .COUT(n26259));
    defparam add_19123_26.INIT0 = 16'h5555;
    defparam add_19123_26.INIT1 = 16'h5555;
    defparam add_19123_26.INJECT1_0 = "NO";
    defparam add_19123_26.INJECT1_1 = "NO";
    CCU2D add_19123_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26257), .COUT(n26258));
    defparam add_19123_24.INIT0 = 16'h5555;
    defparam add_19123_24.INIT1 = 16'h5555;
    defparam add_19123_24.INJECT1_0 = "NO";
    defparam add_19123_24.INJECT1_1 = "NO";
    FD1S3IX count_2618__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i1.GSR = "ENABLED";
    FD1S3IX count_2618__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i2.GSR = "ENABLED";
    FD1S3IX count_2618__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i3.GSR = "ENABLED";
    FD1S3IX count_2618__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i4.GSR = "ENABLED";
    FD1S3IX count_2618__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i5.GSR = "ENABLED";
    FD1S3IX count_2618__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i6.GSR = "ENABLED";
    FD1S3IX count_2618__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i7.GSR = "ENABLED";
    FD1S3IX count_2618__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i8.GSR = "ENABLED";
    FD1S3IX count_2618__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i9.GSR = "ENABLED";
    FD1S3IX count_2618__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i10.GSR = "ENABLED";
    FD1S3IX count_2618__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i11.GSR = "ENABLED";
    FD1S3IX count_2618__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i12.GSR = "ENABLED";
    FD1S3IX count_2618__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i13.GSR = "ENABLED";
    FD1S3IX count_2618__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i14.GSR = "ENABLED";
    FD1S3IX count_2618__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i15.GSR = "ENABLED";
    FD1S3IX count_2618__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i16.GSR = "ENABLED";
    FD1S3IX count_2618__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i17.GSR = "ENABLED";
    FD1S3IX count_2618__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i18.GSR = "ENABLED";
    FD1S3IX count_2618__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i19.GSR = "ENABLED";
    FD1S3IX count_2618__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i20.GSR = "ENABLED";
    FD1S3IX count_2618__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i21.GSR = "ENABLED";
    FD1S3IX count_2618__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i22.GSR = "ENABLED";
    FD1S3IX count_2618__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i23.GSR = "ENABLED";
    FD1S3IX count_2618__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i24.GSR = "ENABLED";
    FD1S3IX count_2618__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i25.GSR = "ENABLED";
    FD1S3IX count_2618__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i26.GSR = "ENABLED";
    FD1S3IX count_2618__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i27.GSR = "ENABLED";
    FD1S3IX count_2618__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i28.GSR = "ENABLED";
    FD1S3IX count_2618__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i29.GSR = "ENABLED";
    FD1S3IX count_2618__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i30.GSR = "ENABLED";
    FD1S3IX count_2618__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16173), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2618__i31.GSR = "ENABLED";
    CCU2D add_19123_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26256), .COUT(n26257));
    defparam add_19123_22.INIT0 = 16'h5555;
    defparam add_19123_22.INIT1 = 16'h5555;
    defparam add_19123_22.INJECT1_0 = "NO";
    defparam add_19123_22.INJECT1_1 = "NO";
    CCU2D add_19123_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26255), .COUT(n26256));
    defparam add_19123_20.INIT0 = 16'h5555;
    defparam add_19123_20.INIT1 = 16'h5555;
    defparam add_19123_20.INJECT1_0 = "NO";
    defparam add_19123_20.INJECT1_1 = "NO";
    CCU2D add_19123_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26254), .COUT(n26255));
    defparam add_19123_18.INIT0 = 16'h5555;
    defparam add_19123_18.INIT1 = 16'h5555;
    defparam add_19123_18.INJECT1_0 = "NO";
    defparam add_19123_18.INJECT1_1 = "NO";
    CCU2D add_19123_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26253), .COUT(n26254));
    defparam add_19123_16.INIT0 = 16'h5555;
    defparam add_19123_16.INIT1 = 16'h5555;
    defparam add_19123_16.INJECT1_0 = "NO";
    defparam add_19123_16.INJECT1_1 = "NO";
    CCU2D add_19123_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26252), .COUT(n26253));
    defparam add_19123_14.INIT0 = 16'h5555;
    defparam add_19123_14.INIT1 = 16'h5555;
    defparam add_19123_14.INJECT1_0 = "NO";
    defparam add_19123_14.INJECT1_1 = "NO";
    CCU2D add_19123_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26251), .COUT(n26252));
    defparam add_19123_12.INIT0 = 16'h5555;
    defparam add_19123_12.INIT1 = 16'h5555;
    defparam add_19123_12.INJECT1_0 = "NO";
    defparam add_19123_12.INJECT1_1 = "NO";
    CCU2D add_19123_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26250), .COUT(n26251));
    defparam add_19123_10.INIT0 = 16'h5aaa;
    defparam add_19123_10.INIT1 = 16'h5555;
    defparam add_19123_10.INJECT1_0 = "NO";
    defparam add_19123_10.INJECT1_1 = "NO";
    CCU2D add_19123_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26249), 
          .COUT(n26250));
    defparam add_19123_8.INIT0 = 16'h5555;
    defparam add_19123_8.INIT1 = 16'h5555;
    defparam add_19123_8.INJECT1_0 = "NO";
    defparam add_19123_8.INJECT1_1 = "NO";
    CCU2D add_19123_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26248), 
          .COUT(n26249));
    defparam add_19123_6.INIT0 = 16'h5aaa;
    defparam add_19123_6.INIT1 = 16'h5aaa;
    defparam add_19123_6.INJECT1_0 = "NO";
    defparam add_19123_6.INJECT1_1 = "NO";
    CCU2D add_19123_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26247), 
          .COUT(n26248));
    defparam add_19123_4.INIT0 = 16'h5555;
    defparam add_19123_4.INIT1 = 16'h5aaa;
    defparam add_19123_4.INJECT1_0 = "NO";
    defparam add_19123_4.INJECT1_1 = "NO";
    CCU2D add_19123_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26247));
    defparam add_19123_2.INIT0 = 16'h1000;
    defparam add_19123_2.INIT1 = 16'h5555;
    defparam add_19123_2.INJECT1_0 = "NO";
    defparam add_19123_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000) 
//

module \ClockDividerP(factor=12000)  (debug_c_c, select_clk, n107, GND_net, 
            n8129, \state[0] , n32380, n30304) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output select_clk;
    input n107;
    input GND_net;
    output n8129;
    input \state[0] ;
    input n32380;
    output n30304;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n34, n24, n38, n32, n2777;
    wire [31:0]n134;
    
    wire n26134, n26133, n26132, n26131, n26130, n26129, n26128, 
        n26127, n26126, n26125, n26124, n26123, n26122, n26121, 
        n26120, n26119, n26231, n26230, n26229, n28703, n26843, 
        n15, n20, n16, n27, n40, n36, n28, n18, n26228, n26227, 
        n26226, n26225, n26224, n26223, n26222, n26221, n26220, 
        n26219;
    
    LUT4 i17_4_lut (.A(count[29]), .B(n34), .C(n24), .D(count[14]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(count[22]), .B(count[21]), .C(count[31]), .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(count[16]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[19]), .B(count[18]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    FD1S3IX count_2617__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2777), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i0.GSR = "ENABLED";
    FD1S3AX clk_o_14 (.D(n107), .CK(debug_c_c), .Q(select_clk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=25, LSE_RCOL=48, LSE_LLINE=21, LSE_RLINE=23 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2617_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26134), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_33.INIT1 = 16'h0000;
    defparam count_2617_add_4_33.INJECT1_0 = "NO";
    defparam count_2617_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26133), .COUT(n26134), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_31.INJECT1_0 = "NO";
    defparam count_2617_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26132), .COUT(n26133), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_29.INJECT1_0 = "NO";
    defparam count_2617_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26131), .COUT(n26132), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_27.INJECT1_0 = "NO";
    defparam count_2617_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26130), .COUT(n26131), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_25.INJECT1_0 = "NO";
    defparam count_2617_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26129), .COUT(n26130), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_23.INJECT1_0 = "NO";
    defparam count_2617_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26128), .COUT(n26129), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_21.INJECT1_0 = "NO";
    defparam count_2617_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26127), .COUT(n26128), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_19.INJECT1_0 = "NO";
    defparam count_2617_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26126), .COUT(n26127), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_17.INJECT1_0 = "NO";
    defparam count_2617_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26125), .COUT(n26126), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_15.INJECT1_0 = "NO";
    defparam count_2617_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26124), .COUT(n26125), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_13.INJECT1_0 = "NO";
    defparam count_2617_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26123), .COUT(n26124), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_11.INJECT1_0 = "NO";
    defparam count_2617_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26122), .COUT(n26123), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_9.INJECT1_0 = "NO";
    defparam count_2617_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26121), .COUT(n26122), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_7.INJECT1_0 = "NO";
    defparam count_2617_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26120), .COUT(n26121), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_5.INJECT1_0 = "NO";
    defparam count_2617_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26119), .COUT(n26120), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2617_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2617_add_4_3.INJECT1_0 = "NO";
    defparam count_2617_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2617_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26119), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617_add_4_1.INIT0 = 16'hF000;
    defparam count_2617_add_4_1.INIT1 = 16'h0555;
    defparam count_2617_add_4_1.INJECT1_0 = "NO";
    defparam count_2617_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_295_4_lut (.A(n8129), .B(select_clk), .C(\state[0] ), 
         .D(n32380), .Z(n30304)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam i1_3_lut_rep_295_4_lut.init = 16'h0002;
    FD1S3IX count_2617__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2777), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i1.GSR = "ENABLED";
    FD1S3IX count_2617__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2777), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i2.GSR = "ENABLED";
    FD1S3IX count_2617__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2777), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i3.GSR = "ENABLED";
    FD1S3IX count_2617__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2777), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i4.GSR = "ENABLED";
    FD1S3IX count_2617__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2777), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i5.GSR = "ENABLED";
    FD1S3IX count_2617__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2777), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i6.GSR = "ENABLED";
    FD1S3IX count_2617__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2777), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i7.GSR = "ENABLED";
    FD1S3IX count_2617__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2777), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i8.GSR = "ENABLED";
    FD1S3IX count_2617__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2777), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i9.GSR = "ENABLED";
    FD1S3IX count_2617__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i10.GSR = "ENABLED";
    FD1S3IX count_2617__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i11.GSR = "ENABLED";
    FD1S3IX count_2617__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i12.GSR = "ENABLED";
    FD1S3IX count_2617__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i13.GSR = "ENABLED";
    FD1S3IX count_2617__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i14.GSR = "ENABLED";
    FD1S3IX count_2617__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i15.GSR = "ENABLED";
    FD1S3IX count_2617__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i16.GSR = "ENABLED";
    FD1S3IX count_2617__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i17.GSR = "ENABLED";
    FD1S3IX count_2617__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i18.GSR = "ENABLED";
    FD1S3IX count_2617__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i19.GSR = "ENABLED";
    FD1S3IX count_2617__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i20.GSR = "ENABLED";
    FD1S3IX count_2617__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i21.GSR = "ENABLED";
    FD1S3IX count_2617__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i22.GSR = "ENABLED";
    FD1S3IX count_2617__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i23.GSR = "ENABLED";
    FD1S3IX count_2617__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i24.GSR = "ENABLED";
    FD1S3IX count_2617__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i25.GSR = "ENABLED";
    FD1S3IX count_2617__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i26.GSR = "ENABLED";
    FD1S3IX count_2617__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i27.GSR = "ENABLED";
    FD1S3IX count_2617__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i28.GSR = "ENABLED";
    FD1S3IX count_2617__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i29.GSR = "ENABLED";
    FD1S3IX count_2617__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i30.GSR = "ENABLED";
    FD1S3IX count_2617__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2777), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2617__i31.GSR = "ENABLED";
    CCU2D add_19122_28 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26231), 
          .S1(n8129));
    defparam add_19122_28.INIT0 = 16'h5555;
    defparam add_19122_28.INIT1 = 16'h0000;
    defparam add_19122_28.INJECT1_0 = "NO";
    defparam add_19122_28.INJECT1_1 = "NO";
    CCU2D add_19122_26 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26230), .COUT(n26231));
    defparam add_19122_26.INIT0 = 16'h5555;
    defparam add_19122_26.INIT1 = 16'h5555;
    defparam add_19122_26.INJECT1_0 = "NO";
    defparam add_19122_26.INJECT1_1 = "NO";
    CCU2D add_19122_24 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26229), .COUT(n26230));
    defparam add_19122_24.INIT0 = 16'h5555;
    defparam add_19122_24.INIT1 = 16'h5555;
    defparam add_19122_24.INJECT1_0 = "NO";
    defparam add_19122_24.INJECT1_1 = "NO";
    LUT4 i21653_2_lut (.A(n28703), .B(n32380), .Z(n2777)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21653_2_lut.init = 16'heeee;
    LUT4 i21651_4_lut (.A(n26843), .B(n15), .C(n20), .D(n16), .Z(n28703)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i21651_4_lut.init = 16'h4000;
    LUT4 i20_4_lut (.A(n27), .B(n40), .C(n36), .D(n28), .Z(n26843)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[11]), .B(count[10]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(count[9]), .B(n18), .C(count[6]), .D(count[7]), 
         .Z(n20)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(count[1]), .B(count[4]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i6_2_lut (.A(count[28]), .B(count[12]), .Z(n27)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    CCU2D add_19122_22 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26228), .COUT(n26229));
    defparam add_19122_22.INIT0 = 16'h5555;
    defparam add_19122_22.INIT1 = 16'h5555;
    defparam add_19122_22.INJECT1_0 = "NO";
    defparam add_19122_22.INJECT1_1 = "NO";
    CCU2D add_19122_20 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26227), .COUT(n26228));
    defparam add_19122_20.INIT0 = 16'h5555;
    defparam add_19122_20.INIT1 = 16'h5555;
    defparam add_19122_20.INJECT1_0 = "NO";
    defparam add_19122_20.INJECT1_1 = "NO";
    CCU2D add_19122_18 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26226), .COUT(n26227));
    defparam add_19122_18.INIT0 = 16'h5555;
    defparam add_19122_18.INIT1 = 16'h5555;
    defparam add_19122_18.INJECT1_0 = "NO";
    defparam add_19122_18.INJECT1_1 = "NO";
    LUT4 i19_4_lut (.A(count[5]), .B(n38), .C(n32), .D(count[20]), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(count[8]), .B(count[25]), .C(count[15]), .D(count[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_4_lut.init = 16'hfffe;
    CCU2D add_19122_16 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26225), .COUT(n26226));
    defparam add_19122_16.INIT0 = 16'h5555;
    defparam add_19122_16.INIT1 = 16'h5555;
    defparam add_19122_16.INJECT1_0 = "NO";
    defparam add_19122_16.INJECT1_1 = "NO";
    LUT4 i7_2_lut (.A(count[17]), .B(count[24]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    CCU2D add_19122_14 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26224), .COUT(n26225));
    defparam add_19122_14.INIT0 = 16'h5555;
    defparam add_19122_14.INIT1 = 16'h5555;
    defparam add_19122_14.INJECT1_0 = "NO";
    defparam add_19122_14.INJECT1_1 = "NO";
    LUT4 i7_4_lut (.A(count[13]), .B(count[2]), .C(count[3]), .D(count[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    CCU2D add_19122_12 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26223), .COUT(n26224));
    defparam add_19122_12.INIT0 = 16'h5555;
    defparam add_19122_12.INIT1 = 16'h5555;
    defparam add_19122_12.INJECT1_0 = "NO";
    defparam add_19122_12.INJECT1_1 = "NO";
    CCU2D add_19122_10 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26222), .COUT(n26223));
    defparam add_19122_10.INIT0 = 16'h5555;
    defparam add_19122_10.INIT1 = 16'h5555;
    defparam add_19122_10.INJECT1_0 = "NO";
    defparam add_19122_10.INJECT1_1 = "NO";
    CCU2D add_19122_8 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26221), .COUT(n26222));
    defparam add_19122_8.INIT0 = 16'h5555;
    defparam add_19122_8.INIT1 = 16'h5aaa;
    defparam add_19122_8.INJECT1_0 = "NO";
    defparam add_19122_8.INJECT1_1 = "NO";
    CCU2D add_19122_6 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26220), .COUT(n26221));
    defparam add_19122_6.INIT0 = 16'h5aaa;
    defparam add_19122_6.INIT1 = 16'h5aaa;
    defparam add_19122_6.INJECT1_0 = "NO";
    defparam add_19122_6.INJECT1_1 = "NO";
    CCU2D add_19122_4 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26219), 
          .COUT(n26220));
    defparam add_19122_4.INIT0 = 16'h5555;
    defparam add_19122_4.INIT1 = 16'h5aaa;
    defparam add_19122_4.INJECT1_0 = "NO";
    defparam add_19122_4.INJECT1_1 = "NO";
    CCU2D add_19122_2 (.A0(count[5]), .B0(count[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26219));
    defparam add_19122_2.INIT0 = 16'h7000;
    defparam add_19122_2.INIT1 = 16'h5aaa;
    defparam add_19122_2.INJECT1_0 = "NO";
    defparam add_19122_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (register_addr, debug_c_c, databus, 
            debug_c_5, \select[4] , n30491, n30489, n30479, n30391, 
            n30488, n30396, n30398, sendcount, n13574, databus_out, 
            n32377, n32379, prev_select, \read_value[1] , rw, n1, 
            n32380, n2673, \select[7] , \sendcount[3] , \select[3] , 
            \select[2] , \select[1] , debug_c_7, n30383, n3806, n5632, 
            n26671, n32376, n30321, \register[1][0] , n97, \register[1][24] , 
            n49, n1307, n28421, n1313, n1310, \register[1][25] , 
            n47, \register[1][29] , n39, n30316, n3666, debug_c_2, 
            debug_c_3, \register[1][30] , n37, debug_c_4, n30324, 
            n21310, n3989, n30344, n3892, n30422, \register_addr[1] , 
            n30411, n30394, n30413, n30385, n17, n4, \reg_size[2] , 
            n30454, \steps_reg[7] , n19, \control_reg[7] , n1_adj_216, 
            \steps_reg[4] , n17_adj_217, n4_adj_218, \steps_reg[6] , 
            n13, n30373, n30417, n28218, n30317, \steps_reg[5] , 
            n14, \steps_reg[3] , n12, \control_reg[7]_adj_219 , n8263, 
            \control_reg[7]_adj_220 , n8272, \reset_count[14] , \reset_count[13] , 
            \reset_count[12] , n26787, n10643, GND_net, uart_rx_c) /* synthesis syn_module_defined=1 */ ;
    output [7:0]register_addr;
    input debug_c_c;
    input [31:0]databus;
    output debug_c_5;
    output \select[4] ;
    output n30491;
    input n30489;
    input n30479;
    output n30391;
    input n30488;
    output n30396;
    output n30398;
    output [4:0]sendcount;
    input n13574;
    output [31:0]databus_out;
    output n32377;
    output n32379;
    input prev_select;
    input \read_value[1] ;
    output rw;
    output n1;
    input n32380;
    output n2673;
    output \select[7] ;
    output \sendcount[3] ;
    output \select[3] ;
    output \select[2] ;
    output \select[1] ;
    output debug_c_7;
    output n30383;
    output n3806;
    output n5632;
    input n26671;
    input n32376;
    input n30321;
    input \register[1][0] ;
    output n97;
    input \register[1][24] ;
    output n49;
    output n1307;
    input n28421;
    output n1313;
    output n1310;
    input \register[1][25] ;
    output n47;
    input \register[1][29] ;
    output n39;
    input n30316;
    output n3666;
    output debug_c_2;
    output debug_c_3;
    input \register[1][30] ;
    output n37;
    output debug_c_4;
    input n30324;
    input n21310;
    output n3989;
    input n30344;
    output n3892;
    output n30422;
    output \register_addr[1] ;
    output n30411;
    output n30394;
    output n30413;
    output n30385;
    input n17;
    input n4;
    input \reg_size[2] ;
    input n30454;
    input \steps_reg[7] ;
    output n19;
    input \control_reg[7] ;
    output n1_adj_216;
    input \steps_reg[4] ;
    output n17_adj_217;
    output n4_adj_218;
    input \steps_reg[6] ;
    output n13;
    input n30373;
    input n30417;
    input n28218;
    output n30317;
    input \steps_reg[5] ;
    output n14;
    input \steps_reg[3] ;
    output n12;
    input \control_reg[7]_adj_219 ;
    output n8263;
    input \control_reg[7]_adj_220 ;
    output n8272;
    input \reset_count[14] ;
    input \reset_count[13] ;
    input \reset_count[12] ;
    input n26787;
    output n10643;
    input GND_net;
    input uart_rx_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire n32376 /* synthesis nomerge= */ ;
    
    wire n2621;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    wire [31:0]n1295;
    
    wire n15359, n30481;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n11, n5, n28067, n26533, n11_adj_423, n11_adj_424, n11_adj_425;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n28329, n11_adj_426;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n11_adj_427, n11_adj_428, n11_adj_429, n11_adj_430, n11_adj_431, 
        n11_adj_432, n11_adj_433, n11_adj_434, n5_adj_435, n28062, 
        n26531, n30486, n10, n30544, n30351, n30402;
    wire [3:0]n1691;
    
    wire n5_adj_436, n28063, n26534, n5_adj_437, n28071, n26647, 
        n30359, n9116, n21586;
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n28330;
    wire [4:0]sendcount_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n30430, n9;
    wire [4:0]n3;
    
    wire n30431, n30400, n5_adj_439, n28069, n26523, n30432;
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n29290, n5_adj_440, n28070, n26648;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n13571;
    wire [7:0]n2037;
    
    wire n30357, n15360;
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    
    wire n29292, n2623, n15974, n1696, n15975, n5_adj_441, n28060, 
        n26502, n5_adj_442, n28072, n26646, n14398, n32388, n27488, 
        n5_adj_443, n28074, n26560, n13277, n5_adj_444, n28073, 
        n26644, n30496, n30495, n30499, n30498, n30318, n30502, 
        n30375, n28059, n30501, n5_adj_445, n28061, n26673, n30505, 
        n30504, n30508, n30507, n30511, n30510, n26682, n5_adj_446, 
        n28075, n26623, n15963, n28360, n30514, n29286, n15965, 
        n30297, n30298, n16045, n30513, n12917;
    wire [7:0]n5623;
    
    wire n30500, n30434, n28589, n21219, n30545, n22, n30517, 
        n5_adj_447, n28057, n26583, n29705, n29706, n30435, n13_adj_448, 
        n27954, escape, n30436, n5_adj_449, n28076, n26641, n30516, 
        n5_adj_450, n28077, n26639, n30520, n30519, n29729, n30542, 
        n30543, n30523, n30522, n30437, n7, n5_adj_452, n28078, 
        n26614, n5_adj_453, n28079, n26637, n5_adj_454, n28080, 
        n26619, n5_adj_455, n28081, n26622, n10550, n5_adj_456, 
        n28082, n26611, n28359, n5_adj_457, n28083, n26640, n5_adj_458, 
        n28084, n26632, n5_adj_459, n28085, n26576, n5_adj_460, 
        n28086, n26579, n5_adj_461, n28088, n26593, n5_adj_462, 
        n28058, n26608, n5_adj_463, n28087, n26600, n30, n28278, 
        n16044, n26676, n1748, n30420, n13012, n8, n27778, n15962, 
        n28310, n15, n15964, n28311, n28032, n28254, n28002, n27666, 
        n28506, n29291, n12888, n11905, n2, n28005, n15968, n15966, 
        send, n2046, busy, n1406, n1407, n11907, n9291, n29902, 
        n1416, n26588, n30524;
    wire [7:0]n9241;
    
    wire n4_c, n9_adj_464, n8_adj_465, n30480, n29901, n30492, n27960, 
        n10_adj_466, n30487, n10747, n12021, n4_adj_467, n4_adj_468, 
        n30426, n6, n28068, n28065, n12_c, n14_c, n27490, n28318, 
        n27630, n27494, n27572, n27506, n27512, n27508, n11_adj_469, 
        n27580, n28476, n9055, n11_adj_470, n27576, n28097;
    wire [7:0]register_addr_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire n11_adj_471, n27628, n27504, n27510, n27574, n27464, n4_adj_472, 
        n30503, n27586, n4_adj_473, n30506, n4_adj_474, n30509, 
        n5_adj_475, n28064, n26538, n4_adj_476, n30515, n5_adj_477, 
        n28066, n26541, n30521, n30518, n30512, n1400, n5_adj_478, 
        n26525, n28232, n5_adj_479, n26535, n5_adj_480, n26529;
    wire [3:0]n9297;
    
    wire n16120, n10768, n18556, n6_adj_481, n5_adj_482, n30493, 
        n30497;
    
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2621), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    LUT4 i14421_2_lut (.A(bufcount[0]), .B(n1295[0]), .Z(n15359)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14421_2_lut.init = 16'h2222;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n30481), .C(\buffer[1] [3]), 
         .D(rx_data[3]), .Z(n11)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2_4_lut (.A(databus[5]), .B(n5), .C(n1295[13]), .D(n28067), 
         .Z(n26533)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 i24_3_lut_4_lut_adj_233 (.A(bufcount[0]), .B(n30481), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_423)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_233.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_234 (.A(bufcount[0]), .B(n30481), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_424)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_234.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_235 (.A(bufcount[0]), .B(n30481), .C(\buffer[1] [6]), 
         .D(rx_data[6]), .Z(n11_adj_425)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_235.init = 16'hf2d0;
    LUT4 select_2088_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1295[4]), 
         .C(rx_data[5]), .D(n28329), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 i24_3_lut_4_lut_adj_236 (.A(bufcount[0]), .B(n30481), .C(rx_data[7]), 
         .D(\buffer[1] [7]), .Z(n11_adj_426)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_236.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_237 (.A(bufcount[0]), .B(n30481), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_adj_427)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_237.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_238 (.A(bufcount[0]), .B(n30481), .C(\buffer[0] [1]), 
         .D(rx_data[1]), .Z(n11_adj_428)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_238.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_239 (.A(bufcount[0]), .B(n30481), .C(rx_data[2]), 
         .D(\buffer[0] [2]), .Z(n11_adj_429)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_239.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_240 (.A(bufcount[0]), .B(n30481), .C(\buffer[0] [3]), 
         .D(rx_data[3]), .Z(n11_adj_430)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_240.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_241 (.A(bufcount[0]), .B(n30481), .C(rx_data[4]), 
         .D(\buffer[0] [4]), .Z(n11_adj_431)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_241.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_242 (.A(bufcount[0]), .B(n30481), .C(\buffer[0] [5]), 
         .D(rx_data[5]), .Z(n11_adj_432)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_242.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_243 (.A(bufcount[0]), .B(n30481), .C(rx_data[6]), 
         .D(\buffer[0] [6]), .Z(n11_adj_433)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_243.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_244 (.A(bufcount[0]), .B(n30481), .C(\buffer[0] [7]), 
         .D(rx_data[7]), .Z(n11_adj_434)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_244.init = 16'hf1e0;
    LUT4 i2_4_lut_adj_245 (.A(databus[6]), .B(n5_adj_435), .C(n1295[13]), 
         .D(n28062), .Z(n26531)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_245.init = 16'hffec;
    LUT4 select_2088_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1295[4]), 
         .C(rx_data[6]), .D(n28329), .Z(n5_adj_435)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 i5_3_lut_4_lut (.A(n30486), .B(n1295[12]), .C(n10), .D(n1295[10]), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_3_lut_4_lut.init = 16'hfffe;
    LUT4 n30375_bdd_4_lut (.A(bufcount[1]), .B(n1295[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n30544)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n30375_bdd_4_lut.init = 16'h0080;
    LUT4 i3285_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n30351), .C(n30402), 
         .D(bufcount[0]), .Z(n1691[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3285_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    LUT4 i2_4_lut_adj_246 (.A(databus[7]), .B(n5_adj_436), .C(n1295[13]), 
         .D(n28063), .Z(n26534)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_246.init = 16'hffec;
    LUT4 select_2088_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1295[4]), 
         .C(rx_data[7]), .D(n28329), .Z(n5_adj_436)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_382_4_lut (.A(\select[4] ), .B(n30491), .C(n30489), 
         .D(n30479), .Z(n30391)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_382_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_387_4_lut (.A(\select[4] ), .B(n30491), .C(n30489), 
         .D(n30488), .Z(n30396)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_387_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_389_4_lut (.A(\select[4] ), .B(n30491), .C(n30489), 
         .D(register_addr[4]), .Z(n30398)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_389_4_lut.init = 16'h0200;
    LUT4 i2_4_lut_adj_247 (.A(databus[8]), .B(n5_adj_437), .C(n1295[13]), 
         .D(n28071), .Z(n26647)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_247.init = 16'hffec;
    FD1P3IX sendcount__i0 (.D(n21586), .SP(n30359), .CD(n9116), .CK(debug_c_c), 
            .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    LUT4 select_2088_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1295[4]), 
         .C(rx_data[0]), .D(n28330), .Z(n5_adj_437)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 i3539_2_lut_rep_421 (.A(sendcount_c[1]), .B(sendcount[0]), .Z(n30430)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3539_2_lut_rep_421.init = 16'h8888;
    LUT4 i14579_3_lut_4_lut (.A(sendcount_c[1]), .B(sendcount[0]), .C(n9), 
         .D(sendcount_c[2]), .Z(n3[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;
    defparam i14579_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i3542_2_lut_rep_422 (.A(sendcount_c[1]), .B(sendcount[0]), .Z(n30431)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3542_2_lut_rep_422.init = 16'heeee;
    LUT4 i1_2_lut_rep_391_3_lut (.A(sendcount_c[1]), .B(sendcount[0]), .C(sendcount_c[2]), 
         .Z(n30400)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_391_3_lut.init = 16'h1e1e;
    LUT4 i2_4_lut_adj_248 (.A(databus[9]), .B(n5_adj_439), .C(n1295[13]), 
         .D(n28069), .Z(n26523)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_248.init = 16'hffec;
    LUT4 i3329_2_lut_rep_423 (.A(sendcount_c[1]), .B(sendcount[0]), .Z(n30432)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i3329_2_lut_rep_423.init = 16'h9999;
    LUT4 select_2088_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1295[4]), 
         .C(rx_data[1]), .D(n28330), .Z(n5_adj_439)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i14580_2_lut_2_lut_3_lut (.A(sendcount_c[1]), .B(sendcount[0]), 
         .C(n9), .Z(n3[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i14580_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 n12668_bdd_4_lut_22043_4_lut (.A(sendcount_c[1]), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n29290)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n12668_bdd_4_lut_22043_4_lut.init = 16'h6420;
    LUT4 i2_4_lut_adj_249 (.A(databus[10]), .B(n5_adj_440), .C(n1295[13]), 
         .D(n28070), .Z(n26648)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_249.init = 16'hffec;
    LUT4 select_2088_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1295[4]), 
         .C(rx_data[2]), .D(n28330), .Z(n5_adj_440)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_26_i5_4_lut.init = 16'h88c0;
    FD1P3AX tx_data_i0_i0 (.D(n2037[0]), .SP(n13571), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n15360), .CK(debug_c_c), .CD(n30357), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n29292), .SP(n13574), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    PFUMX i9563 (.BLUT(n15974), .ALUT(n1691[1]), .C0(n1696), .Z(n15975));
    LUT4 i2_4_lut_adj_250 (.A(databus[11]), .B(n5_adj_441), .C(n1295[13]), 
         .D(n28060), .Z(n26502)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_250.init = 16'hffec;
    LUT4 select_2088_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1295[4]), 
         .C(rx_data[3]), .D(n28330), .Z(n5_adj_441)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_251 (.A(databus[12]), .B(n5_adj_442), .C(n1295[13]), 
         .D(n28072), .Z(n26646)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_251.init = 16'hffec;
    LUT4 select_2088_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1295[4]), 
         .C(rx_data[4]), .D(n28330), .Z(n5_adj_442)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_28_i5_4_lut.init = 16'h88c0;
    FD1P3IX buffer_0___i1 (.D(n27488), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_252 (.A(databus[13]), .B(n5_adj_443), .C(n1295[13]), 
         .D(n28074), .Z(n26560)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_252.init = 16'hffec;
    FD1S3JX state_FSM_i1 (.D(n13277), .CK(debug_c_c), .PD(n32388), .Q(n1295[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 select_2088_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1295[4]), 
         .C(rx_data[5]), .D(n28330), .Z(n5_adj_443)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_253 (.A(databus[14]), .B(n5_adj_444), .C(n1295[13]), 
         .D(n28073), .Z(n26644)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_253.init = 16'hffec;
    LUT4 i1_4_lut_then_4_lut (.A(esc_data[6]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[4]), .Z(n30496)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0400;
    LUT4 i1_4_lut_else_4_lut (.A(esc_data[6]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[4]), .Z(n30495)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 select_2088_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1295[4]), 
         .C(rx_data[6]), .D(n28330), .Z(n5_adj_444)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i9559_then_4_lut (.A(bufcount[3]), .B(n1295[0]), .C(n1295[3]), 
         .D(n1295[4]), .Z(n30499)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i9559_then_4_lut.init = 16'haaa2;
    LUT4 i9559_else_4_lut (.A(bufcount[3]), .B(n1295[0]), .C(n1295[3]), 
         .D(n1295[4]), .Z(n30498)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i9559_else_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_309_3_lut_4_lut (.A(n32377), .B(n30398), .C(n32379), 
         .D(prev_select), .Z(n30318)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_309_3_lut_4_lut.init = 16'h0008;
    LUT4 i14886_2_lut (.A(bufcount[1]), .B(n1295[0]), .Z(n15974)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14886_2_lut.init = 16'h2222;
    LUT4 i21459_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(sendcount_c[1]), 
         .Z(n30502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21459_then_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut (.A(n1295[3]), .B(n30375), .C(\buffer[2] [2]), 
         .Z(n28059)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i21459_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(sendcount_c[1]), 
         .Z(n30501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21459_else_3_lut.init = 16'hcaca;
    LUT4 Select_4226_i1_2_lut_3_lut_4_lut (.A(n32377), .B(n30398), .C(\read_value[1] ), 
         .D(rw), .Z(n1)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4226_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_254 (.A(databus[15]), .B(n5_adj_445), .C(n1295[13]), 
         .D(n28061), .Z(n26673)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_254.init = 16'hffec;
    LUT4 i21462_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(sendcount_c[1]), 
         .Z(n30505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21462_then_3_lut.init = 16'hcaca;
    LUT4 i21462_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(sendcount_c[1]), 
         .Z(n30504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21462_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n30398), .C(n32380), 
         .D(prev_select), .Z(n2673)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 select_2088_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1295[4]), 
         .C(rx_data[7]), .D(n28330), .Z(n5_adj_445)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i21465_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(sendcount_c[1]), 
         .Z(n30508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21465_then_3_lut.init = 16'hcaca;
    LUT4 i21465_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(sendcount_c[1]), 
         .Z(n30507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21465_else_3_lut.init = 16'hcaca;
    LUT4 i21468_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(sendcount_c[1]), 
         .Z(n30511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21468_then_3_lut.init = 16'hcaca;
    LUT4 i21468_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(sendcount_c[1]), 
         .Z(n30510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21468_else_3_lut.init = 16'hcaca;
    PFUMX i8948 (.BLUT(n15359), .ALUT(n26682), .C0(n1696), .Z(n15360));
    LUT4 i2_4_lut_adj_255 (.A(databus[16]), .B(n5_adj_446), .C(n1295[13]), 
         .D(n28075), .Z(n26623)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_255.init = 16'hffec;
    FD1S3IX select__i7 (.D(n15963), .CK(debug_c_c), .CD(n32388), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 select_2088_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1295[4]), 
         .C(rx_data[0]), .D(n28360), .Z(n5_adj_446)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 i21471_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(sendcount_c[1]), 
         .Z(n30514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21471_then_3_lut.init = 16'hcaca;
    LUT4 n12668_bdd_2_lut_22039 (.A(sendcount[0]), .B(\sendcount[3] ), .Z(n29286)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n12668_bdd_2_lut_22039.init = 16'hbbbb;
    FD1S3IX select__i4 (.D(n15965), .CK(debug_c_c), .CD(n32388), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1S3IX select__i3 (.D(n30297), .CK(debug_c_c), .CD(n32388), .Q(\select[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i3.GSR = "ENABLED";
    FD1S3IX select__i2 (.D(n30298), .CK(debug_c_c), .CD(n32388), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1S3IX select__i1 (.D(n16045), .CK(debug_c_c), .CD(n32388), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    LUT4 i21471_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(sendcount_c[1]), 
         .Z(n30513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21471_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_256 (.A(rx_data[1]), .B(rx_data[4]), .C(rx_data[3]), 
         .Z(n12917)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_3_lut_adj_256.init = 16'h0808;
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2623), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i4 (.D(n5623[4]), .SP(n13574), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n5623[2]), .SP(n13574), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n5623[1]), .SP(n13574), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    FD1S3IX bufcount__i3 (.D(n30500), .CK(debug_c_c), .CD(n32388), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    LUT4 i21302_2_lut_rep_425 (.A(rx_data[7]), .B(rx_data[6]), .Z(n30434)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21302_2_lut_rep_425.init = 16'heeee;
    LUT4 i21448_3_lut_rep_366_4_lut (.A(rx_data[7]), .B(rx_data[6]), .C(n28589), 
         .D(n21219), .Z(n30375)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21448_3_lut_rep_366_4_lut.init = 16'hfffe;
    FD1S3IX bufcount__i2 (.D(n30545), .CK(debug_c_c), .CD(n32388), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n15975), .CK(debug_c_c), .CD(n32388), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2037[4]), .SP(n13571), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n22), .SP(n13571), .CK(debug_c_c), .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2037[1]), .SP(n13571), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    LUT4 i21474_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(sendcount_c[1]), 
         .Z(n30517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21474_then_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_257 (.A(databus[17]), .B(n5_adj_447), .C(n1295[13]), 
         .D(n28057), .Z(n26583)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_257.init = 16'hffec;
    LUT4 sendcount_4__bdd_3_lut (.A(sendcount_c[4]), .B(n29705), .C(\sendcount[3] ), 
         .Z(n29706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut.init = 16'hcaca;
    LUT4 select_2088_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1295[4]), 
         .C(rx_data[1]), .D(n28360), .Z(n5_adj_447)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_426 (.A(rx_data[5]), .B(rx_data[0]), .Z(n30435)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i1_2_lut_rep_426.init = 16'hbbbb;
    LUT4 i2_3_lut_4_lut (.A(rx_data[5]), .B(rx_data[0]), .C(rx_data[2]), 
         .D(n13_adj_448), .Z(n27954)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i2_3_lut_4_lut.init = 16'hfffb;
    LUT4 i907_2_lut_rep_427 (.A(escape), .B(debug_c_7), .Z(n30436)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i907_2_lut_rep_427.init = 16'hbbbb;
    LUT4 i2_4_lut_adj_258 (.A(databus[18]), .B(n5_adj_449), .C(n1295[13]), 
         .D(n28076), .Z(n26641)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_258.init = 16'hffec;
    LUT4 select_2088_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1295[4]), 
         .C(rx_data[2]), .D(n28360), .Z(n5_adj_449)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 i21474_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(sendcount_c[1]), 
         .Z(n30516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21474_else_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_259 (.A(databus[19]), .B(n5_adj_450), .C(n1295[13]), 
         .D(n28077), .Z(n26639)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_259.init = 16'hffec;
    LUT4 sendcount_4__bdd_4_lut (.A(sendcount_c[4]), .B(sendcount_c[2]), 
         .C(sendcount_c[1]), .D(sendcount[0]), .Z(n29705)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_4__bdd_4_lut.init = 16'h6aaa;
    LUT4 i938_3_lut (.A(n1295[5]), .B(n30383), .C(n1295[10]), .Z(n2621)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i938_3_lut.init = 16'hc8c8;
    LUT4 select_2088_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1295[4]), 
         .C(rx_data[3]), .D(n28360), .Z(n5_adj_450)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 i21477_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(sendcount_c[1]), 
         .Z(n30520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21477_then_3_lut.init = 16'hcaca;
    LUT4 i21477_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(sendcount_c[1]), 
         .Z(n30519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21477_else_3_lut.init = 16'hcaca;
    LUT4 rx_data_3__bdd_4_lut_22702 (.A(rx_data[3]), .B(rx_data[2]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n29729)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_3__bdd_4_lut_22702.init = 16'h6001;
    FD1P3IX sendcount__i4 (.D(n29706), .SP(n30359), .CD(n9116), .CK(debug_c_c), 
            .Q(sendcount_c[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 n30542_bdd_2_lut (.A(n30542), .B(n1295[4]), .Z(n30543)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n30542_bdd_2_lut.init = 16'heeee;
    LUT4 n30375_bdd_4_lut_22357 (.A(n30375), .B(n30436), .C(n1295[0]), 
         .D(n1295[3]), .Z(n30542)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n30375_bdd_4_lut_22357.init = 16'hee0f;
    LUT4 i21948_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(sendcount_c[1]), 
         .Z(n30523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21948_then_3_lut.init = 16'hcaca;
    LUT4 i21948_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(sendcount_c[1]), 
         .Z(n30522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21948_else_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_342_4_lut (.A(escape), .B(debug_c_7), .C(n30375), 
         .D(n1295[4]), .Z(n30351)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_342_4_lut.init = 16'hfffb;
    FD1P3IX sendcount__i3 (.D(n3[3]), .SP(n30359), .CD(n9116), .CK(debug_c_c), 
            .Q(\sendcount[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3IX sendcount__i2 (.D(n3[2]), .SP(n30359), .CD(n9116), .CK(debug_c_c), 
            .Q(sendcount_c[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n3[1]), .SP(n30359), .CD(n9116), .CK(debug_c_c), 
            .Q(sendcount_c[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 i1_3_lut_rep_428 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n30437)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_rep_428.init = 16'hecec;
    LUT4 i2_2_lut_rep_393_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1295[4]), .Z(n30402)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_393_4_lut.init = 16'hecff;
    LUT4 i1_2_lut_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1295[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hec00;
    LUT4 i2_4_lut_adj_260 (.A(databus[20]), .B(n5_adj_452), .C(n1295[13]), 
         .D(n28078), .Z(n26614)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_260.init = 16'hffec;
    LUT4 select_2088_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1295[4]), 
         .C(rx_data[4]), .D(n28360), .Z(n5_adj_452)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_261 (.A(databus[21]), .B(n5_adj_453), .C(n1295[13]), 
         .D(n28079), .Z(n26637)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_261.init = 16'hffec;
    LUT4 select_2088_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1295[4]), 
         .C(rx_data[5]), .D(n28360), .Z(n5_adj_453)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_262 (.A(databus[22]), .B(n5_adj_454), .C(n1295[13]), 
         .D(n28080), .Z(n26619)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_262.init = 16'hffec;
    LUT4 select_2088_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1295[4]), 
         .C(rx_data[6]), .D(n28360), .Z(n5_adj_454)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_263 (.A(databus[23]), .B(n5_adj_455), .C(n1295[13]), 
         .D(n28081), .Z(n26622)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_263.init = 16'hffec;
    LUT4 select_2088_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1295[4]), 
         .C(rx_data[7]), .D(n28360), .Z(n5_adj_455)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_39_i5_4_lut.init = 16'h88c0;
    FD1S3AX escape_501 (.D(n10550), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_264 (.A(databus[24]), .B(n5_adj_456), .C(n1295[13]), 
         .D(n28082), .Z(n26611)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_264.init = 16'hffec;
    LUT4 select_2088_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1295[4]), 
         .C(rx_data[0]), .D(n28359), .Z(n5_adj_456)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_265 (.A(databus[25]), .B(n5_adj_457), .C(n1295[13]), 
         .D(n28083), .Z(n26640)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_265.init = 16'hffec;
    LUT4 select_2088_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1295[4]), 
         .C(rx_data[1]), .D(n28359), .Z(n5_adj_457)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_41_i5_4_lut.init = 16'h88c0;
    FD1P3AX rw_498 (.D(n1295[10]), .SP(n2621), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_266 (.A(databus[26]), .B(n5_adj_458), .C(n1295[13]), 
         .D(n28084), .Z(n26632)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_266.init = 16'hffec;
    LUT4 select_2088_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1295[4]), 
         .C(rx_data[2]), .D(n28359), .Z(n5_adj_458)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_267 (.A(databus[27]), .B(n5_adj_459), .C(n1295[13]), 
         .D(n28085), .Z(n26576)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_267.init = 16'hffec;
    LUT4 select_2088_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1295[4]), 
         .C(rx_data[3]), .D(n28359), .Z(n5_adj_459)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_268 (.A(databus[28]), .B(n5_adj_460), .C(n1295[13]), 
         .D(n28086), .Z(n26579)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_268.init = 16'hffec;
    LUT4 select_2088_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1295[4]), 
         .C(rx_data[4]), .D(n28359), .Z(n5_adj_460)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_269 (.A(databus[29]), .B(n5_adj_461), .C(n1295[13]), 
         .D(n28088), .Z(n26593)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_269.init = 16'hffec;
    LUT4 select_2088_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1295[4]), 
         .C(rx_data[5]), .D(n28359), .Z(n5_adj_461)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_270 (.A(databus[30]), .B(n5_adj_462), .C(n1295[13]), 
         .D(n28058), .Z(n26608)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_270.init = 16'hffec;
    LUT4 select_2088_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1295[4]), 
         .C(rx_data[6]), .D(n28359), .Z(n5_adj_462)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_271 (.A(databus[31]), .B(n5_adj_463), .C(n1295[13]), 
         .D(n28087), .Z(n26600)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_271.init = 16'hffec;
    LUT4 i2_3_lut_4_lut_adj_272 (.A(register_addr[5]), .B(n30), .C(n30318), 
         .D(n28278), .Z(n3806)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_272.init = 16'h8000;
    LUT4 select_2088_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1295[4]), 
         .C(rx_data[7]), .D(n28359), .Z(n5_adj_463)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_47_i5_4_lut.init = 16'h88c0;
    PFUMX i9633 (.BLUT(n16044), .ALUT(n26676), .C0(n1748), .Z(n16045));
    LUT4 i1_4_lut (.A(n30420), .B(debug_c_7), .C(n13012), .D(n8), .Z(n27778)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'hdc50;
    PFUMX i9551 (.BLUT(n15962), .ALUT(n28310), .C0(n1748), .Z(n15963));
    LUT4 i1_3_lut (.A(n15), .B(n1295[1]), .C(n1295[0]), .Z(n8)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    PFUMX i9553 (.BLUT(n15964), .ALUT(n28311), .C0(n1748), .Z(n15965));
    LUT4 i3_4_lut (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), .D(n27954), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_273 (.A(n1295[3]), .B(n28032), .C(rx_data[2]), .D(n28254), 
         .Z(n13012)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3_4_lut_adj_273.init = 16'h8000;
    LUT4 i2_4_lut_adj_274 (.A(escape), .B(n13_adj_448), .C(debug_c_7), 
         .D(n12917), .Z(n28032)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2_4_lut_adj_274.init = 16'h1000;
    LUT4 i1_2_lut (.A(rx_data[0]), .B(rx_data[5]), .Z(n28254)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_275 (.A(n1295[4]), .B(debug_c_7), .C(n1295[2]), 
         .D(n28002), .Z(n27666)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_275.init = 16'heeea;
    LUT4 i1_4_lut_adj_276 (.A(n15), .B(n1295[3]), .C(n1295[0]), .D(n28506), 
         .Z(n28002)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_276.init = 16'h50dc;
    PFUMX i21950 (.BLUT(n29291), .ALUT(n29286), .C0(n5632), .Z(n29292));
    LUT4 i21358_3_lut (.A(n12888), .B(escape), .C(n15), .Z(n28506)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i21358_3_lut.init = 16'hecec;
    LUT4 i5496_3_lut (.A(debug_c_7), .B(n1295[3]), .C(n1295[2]), .Z(n11905)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5496_3_lut.init = 16'h5454;
    LUT4 i21813_3_lut (.A(debug_c_7), .B(n2), .C(n1295[3]), .Z(n28005)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i21813_3_lut.init = 16'h2020;
    LUT4 i3_4_lut_adj_277 (.A(escape), .B(n30434), .C(n29729), .D(n28254), 
         .Z(n2)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_277.init = 16'h1000;
    LUT4 i14821_2_lut_3_lut (.A(n1295[0]), .B(n1295[8]), .C(\select[1] ), 
         .Z(n16044)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14821_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_278 (.A(n1295[0]), .B(n1295[8]), .C(\select[4] ), 
         .Z(n15964)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_278.init = 16'h1010;
    LUT4 i14894_2_lut_3_lut (.A(n1295[0]), .B(n1295[8]), .C(\select[2] ), 
         .Z(n15968)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14894_2_lut_3_lut.init = 16'h1010;
    LUT4 i14532_2_lut_3_lut (.A(n1295[0]), .B(n1295[8]), .C(\select[7] ), 
         .Z(n15962)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14532_2_lut_3_lut.init = 16'h1010;
    LUT4 i14424_2_lut_3_lut (.A(n1295[0]), .B(n1295[8]), .C(\select[3] ), 
         .Z(n15966)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14424_2_lut_3_lut.init = 16'h1010;
    FD1P3IX send_491 (.D(n32376), .SP(n2046), .CD(n26671), .CK(debug_c_c), 
            .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_279 (.A(register_addr[0]), .B(n30321), .C(\register[1][0] ), 
         .Z(n97)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_279.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_280 (.A(register_addr[0]), .B(n30321), .C(\register[1][24] ), 
         .Z(n49)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_280.init = 16'h2020;
    LUT4 i1_2_lut_adj_281 (.A(register_addr[4]), .B(register_addr[3]), .Z(n28278)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_281.init = 16'h2222;
    LUT4 reduce_or_457_i1_3_lut (.A(busy), .B(n1295[13]), .C(n1307), .Z(n1406)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_457_i1_3_lut.init = 16'hdcdc;
    LUT4 i3_4_lut_adj_282 (.A(register_addr[2]), .B(n30491), .C(n32380), 
         .D(n28421), .Z(n30)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_adj_282.init = 16'h0100;
    LUT4 i459_2_lut (.A(n5632), .B(n1313), .Z(n1407)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i459_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_283 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n28360)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_283.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_284 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n28359)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_284.init = 16'hbfbf;
    LUT4 i5497_3_lut (.A(busy), .B(n1310), .C(n1295[16]), .Z(n11907)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5497_3_lut.init = 16'ha8a8;
    LUT4 i2_4_lut_adj_285 (.A(n9291), .B(n29902), .C(n1295[15]), .D(n1416), 
         .Z(n26588)) /* synthesis lut_function=(A (B+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_285.init = 16'hffdc;
    LUT4 n29290_bdd_3_lut_4_lut (.A(sendcount_c[2]), .B(n30431), .C(n30524), 
         .D(n29290), .Z(n29291)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n29290_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 i1_2_lut_3_lut_adj_286 (.A(register_addr[0]), .B(n30321), .C(\register[1][25] ), 
         .Z(n47)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_286.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_287 (.A(register_addr[0]), .B(n30321), .C(\register[1][29] ), 
         .Z(n39)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_287.init = 16'h2020;
    LUT4 i2_3_lut_4_lut_adj_288 (.A(n32377), .B(n30), .C(n30316), .D(n28278), 
         .Z(n3666)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_288.init = 16'h4000;
    LUT4 i468_2_lut (.A(busy), .B(n1310), .Z(n1416)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i468_2_lut.init = 16'h4444;
    LUT4 mux_1861_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n5632), 
         .Z(n5623[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1861_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_c)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 i5_4_lut (.A(n9_adj_464), .B(n1295[15]), .C(n8_adj_465), .D(n1295[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_289 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n28329)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_289.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_290 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n28330)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_290.init = 16'hbfbf;
    LUT4 i2_2_lut (.A(n1295[9]), .B(n1310), .Z(n8_adj_465)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_471 (.A(n1313), .B(sendcount_c[4]), .Z(n30480)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_471.init = 16'h2222;
    LUT4 motor_pwm_r_c_bdd_2_lut_22157_3_lut (.A(n1313), .B(sendcount_c[4]), 
         .C(n29901), .Z(n29902)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam motor_pwm_r_c_bdd_2_lut_22157_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_else_4_lut_adj_291 (.A(sendcount_c[4]), .B(sendcount[0]), 
         .C(sendcount_c[1]), .D(sendcount_c[2]), .Z(n30492)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut_adj_291.init = 16'h4001;
    LUT4 i2_3_lut (.A(n1295[13]), .B(n1295[7]), .C(n1295[5]), .Z(n27960)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i3235_2_lut_rep_472 (.A(bufcount[1]), .B(bufcount[2]), .Z(n30481)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3235_2_lut_rep_472.init = 16'heeee;
    LUT4 mux_1861_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n5632), 
         .Z(n5623[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1861_i3_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_292 (.A(n1295[10]), .B(n30486), .C(n10_adj_466), 
         .D(n30487), .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_292.init = 16'hfffe;
    LUT4 i1_3_lut_adj_293 (.A(n1295[18]), .B(n1295[19]), .C(busy), .Z(n10747)) /* synthesis lut_function=(A+!((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_adj_293.init = 16'haeae;
    LUT4 i5610_3_lut (.A(busy), .B(n1307), .C(n1295[19]), .Z(n12021)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5610_3_lut.init = 16'ha8a8;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_467)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i2870_2_lut_rep_411_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n30420)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2870_2_lut_rep_411_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_294 (.A(register_addr[0]), .B(n30321), .C(\register[1][30] ), 
         .Z(n37)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_294.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1295[4]), .B(n30437), .C(bufcount[0]), 
         .D(n30351), .Z(n26682)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hd222;
    LUT4 mux_1861_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n5632), 
         .Z(n5623[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1861_i2_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut (.A(n1295[18]), .B(n1295[2]), .C(n1295[6]), .D(n1295[7]), 
         .Z(n10_adj_466)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_adj_468)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 i4_4_lut_adj_295 (.A(n1295[6]), .B(n30426), .C(n27960), .D(n6), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4_4_lut_adj_295.init = 16'hfffe;
    LUT4 i1_2_lut_adj_296 (.A(n1295[4]), .B(n1307), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_296.init = 16'heeee;
    LUT4 i4_4_lut_adj_297 (.A(n1295[11]), .B(n1295[9]), .C(n1295[8]), 
         .D(n1295[13]), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_297.init = 16'hfffe;
    LUT4 i4_2_lut_rep_477 (.A(n1313), .B(n1295[15]), .Z(n30486)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_477.init = 16'heeee;
    LUT4 i1_2_lut_rep_417_3_lut (.A(n1313), .B(n1295[15]), .C(n1295[12]), 
         .Z(n30426)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_417_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_478 (.A(n1295[19]), .B(n1295[3]), .C(n1295[11]), 
         .Z(n30487)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_rep_478.init = 16'hfefe;
    LUT4 i3_2_lut_4_lut (.A(n1295[19]), .B(n1295[3]), .C(n1295[11]), .D(n27960), 
         .Z(n9_adj_464)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_298 (.A(n32377), .B(n30), .C(n30324), .D(n21310), 
         .Z(n3989)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_298.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_adj_299 (.A(n1295[3]), .B(n30375), .C(\buffer[2] [3]), 
         .Z(n28068)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_299.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_300 (.A(n1295[3]), .B(n30375), .C(\buffer[2] [4]), 
         .Z(n28065)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_300.init = 16'h8080;
    LUT4 i21743_3_lut_4_lut (.A(n12_c), .B(\buffer[0] [2]), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n28310)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i21743_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_301 (.A(n1295[4]), .B(\buffer[0] [1]), .C(n11_adj_428), 
         .D(n14_c), .Z(n27490)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_301.init = 16'heca0;
    LUT4 i21754_3_lut_4_lut (.A(n12_c), .B(\buffer[0] [2]), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n28311)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i21754_3_lut_4_lut.init = 16'h0004;
    LUT4 i21712_3_lut_4_lut (.A(\buffer[0] [2]), .B(n12_c), .C(\buffer[0] [0]), 
         .D(\buffer[0] [1]), .Z(n26676)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i21712_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_302 (.A(\buffer[0] [2]), .B(n12_c), .C(\buffer[0] [1]), 
         .Z(n28318)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i1_2_lut_3_lut_adj_302.init = 16'hefef;
    LUT4 i1_4_lut_adj_303 (.A(n1295[4]), .B(\buffer[0] [0]), .C(n11_adj_427), 
         .D(n14_c), .Z(n27488)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_303.init = 16'heca0;
    LUT4 i1_4_lut_adj_304 (.A(n1295[4]), .B(\buffer[0] [2]), .C(n11_adj_429), 
         .D(n14_c), .Z(n27630)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_304.init = 16'heca0;
    LUT4 i1_4_lut_adj_305 (.A(n1295[4]), .B(\buffer[0] [3]), .C(n11_adj_430), 
         .D(n14_c), .Z(n27494)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_305.init = 16'heca0;
    LUT4 i1_4_lut_adj_306 (.A(n1295[4]), .B(\buffer[0] [4]), .C(n11_adj_431), 
         .D(n14_c), .Z(n27572)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_306.init = 16'heca0;
    LUT4 i1_4_lut_adj_307 (.A(n1295[4]), .B(\buffer[0] [5]), .C(n11_adj_432), 
         .D(n14_c), .Z(n27506)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_307.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_adj_308 (.A(n1295[3]), .B(n30375), .C(\buffer[2] [5]), 
         .Z(n28067)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_308.init = 16'h8080;
    LUT4 i1_4_lut_adj_309 (.A(n1295[4]), .B(\buffer[0] [6]), .C(n11_adj_433), 
         .D(n14_c), .Z(n27512)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_309.init = 16'heca0;
    LUT4 i1_4_lut_adj_310 (.A(n1295[4]), .B(\buffer[0] [7]), .C(n11_adj_434), 
         .D(n14_c), .Z(n27508)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_310.init = 16'heca0;
    LUT4 i1_4_lut_adj_311 (.A(n1295[4]), .B(\buffer[1] [0]), .C(n11_adj_469), 
         .D(n14_c), .Z(n27580)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_311.init = 16'heca0;
    LUT4 i21784_4_lut (.A(n7), .B(n28476), .C(n30436), .D(n1295[3]), 
         .Z(n9055)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i21784_4_lut.init = 16'h0544;
    LUT4 i21329_3_lut (.A(n1295[13]), .B(n1295[0]), .C(n1295[4]), .Z(n28476)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i21329_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut_adj_312 (.A(n32377), .B(n30), .C(n30344), .D(n21310), 
         .Z(n3892)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_312.init = 16'h0080;
    LUT4 i1_4_lut_adj_313 (.A(n1295[4]), .B(\buffer[1] [1]), .C(n11_adj_470), 
         .D(n14_c), .Z(n27576)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_313.init = 16'heca0;
    LUT4 i1_4_lut_adj_314 (.A(n28097), .B(debug_c_7), .C(n1295[0]), .D(n1295[1]), 
         .Z(n13277)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_314.init = 16'hbbba;
    LUT4 i1_2_lut_rep_482 (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .Z(n30491)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_482.init = 16'heeee;
    LUT4 i3_4_lut_adj_315 (.A(\sendcount[3] ), .B(n30431), .C(sendcount_c[2]), 
         .D(n30480), .Z(n28097)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_315.init = 16'h0200;
    LUT4 i1_4_lut_adj_316 (.A(n1295[4]), .B(\buffer[1] [2]), .C(n11_adj_471), 
         .D(n14_c), .Z(n27628)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_316.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_adj_317 (.A(n1295[3]), .B(n30375), .C(\buffer[2] [6]), 
         .Z(n28062)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_317.init = 16'h8080;
    LUT4 i1_4_lut_adj_318 (.A(n1295[4]), .B(\buffer[1] [3]), .C(n11), 
         .D(n14_c), .Z(n27504)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_318.init = 16'heca0;
    LUT4 i1_4_lut_adj_319 (.A(n1295[4]), .B(\buffer[1] [4]), .C(n11_adj_423), 
         .D(n14_c), .Z(n27510)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_319.init = 16'heca0;
    LUT4 i1_4_lut_adj_320 (.A(n1295[4]), .B(\buffer[1] [5]), .C(n11_adj_424), 
         .D(n14_c), .Z(n27574)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_320.init = 16'heca0;
    LUT4 i1_4_lut_adj_321 (.A(n1295[4]), .B(\buffer[1] [6]), .C(n11_adj_425), 
         .D(n14_c), .Z(n27464)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_321.init = 16'heca0;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n30432), .B(n30400), .C(n4_adj_472), 
         .D(n30503), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_4_lut_adj_322 (.A(n1295[4]), .B(\buffer[1] [7]), .C(n11_adj_426), 
         .D(n14_c), .Z(n27586)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_322.init = 16'heca0;
    LUT4 i1_2_lut_rep_413_3_lut_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(n32377), .D(register_addr[4]), .Z(n30422)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_413_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_rep_402_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(register_addr[0]), .D(\register_addr[1] ), .Z(n30411)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_rep_402_4_lut.init = 16'h0100;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n30432), .B(n30400), .C(n4_adj_473), 
         .D(n30506), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i21316_2_lut_rep_385_3_lut_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(register_addr[3]), .D(register_addr[5]), .Z(n30394)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i21316_2_lut_rep_385_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n30432), .B(n30400), .C(n4_adj_474), 
         .D(n30509), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i2_4_lut_adj_323 (.A(databus[0]), .B(n5_adj_475), .C(n1295[13]), 
         .D(n28064), .Z(n26538)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_323.init = 16'hffec;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n30432), .B(n30400), .C(n4_adj_476), 
         .D(n30515), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 select_2088_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1295[4]), 
         .C(rx_data[0]), .D(n28329), .Z(n5_adj_475)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 n28096_bdd_4_lut (.A(\sendcount[3] ), .B(sendcount[0]), .C(sendcount_c[1]), 
         .D(sendcount_c[2]), .Z(n29901)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n28096_bdd_4_lut.init = 16'h4001;
    LUT4 i2_4_lut_adj_324 (.A(databus[1]), .B(n5_adj_477), .C(n1295[13]), 
         .D(n28066), .Z(n26541)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_324.init = 16'hffec;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n30432), .B(n30400), .C(n4_adj_468), 
         .D(n30521), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n30432), .B(n30400), .C(n4_adj_467), 
         .D(n30518), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n30432), .B(n30400), .C(n4_c), 
         .D(n30512), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 select_2088_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1295[4]), 
         .C(rx_data[1]), .D(n28329), .Z(n5_adj_477)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i14551_2_lut_rep_404_3_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(n32377), .Z(n30413)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14551_2_lut_rep_404_3_lut.init = 16'hfefe;
    LUT4 reduce_or_451_i1_3_lut_4_lut (.A(n30420), .B(n13012), .C(\buffer[0] [7]), 
         .D(n1295[9]), .Z(n1400)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_451_i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i4527_2_lut_rep_376_3_lut_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(register_addr[4]), .D(n32377), .Z(n30385)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4527_2_lut_rep_376_3_lut_4_lut.init = 16'h0010;
    LUT4 i2_4_lut_adj_325 (.A(databus[2]), .B(n5_adj_478), .C(n1295[13]), 
         .D(n28059), .Z(n26525)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_325.init = 16'hffec;
    LUT4 select_2088_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1295[4]), 
         .C(rx_data[2]), .D(n28329), .Z(n5_adj_478)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n30481), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n13012), .Z(n28232)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i2_4_lut_adj_326 (.A(databus[3]), .B(n5_adj_479), .C(n1295[13]), 
         .D(n28068), .Z(n26535)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_326.init = 16'hffec;
    LUT4 select_2088_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1295[4]), 
         .C(rx_data[3]), .D(n28329), .Z(n5_adj_479)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_327 (.A(databus[4]), .B(n5_adj_480), .C(n1295[13]), 
         .D(n28065), .Z(n26529)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_327.init = 16'hffec;
    LUT4 select_2088_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1295[4]), 
         .C(rx_data[4]), .D(n28329), .Z(n5_adj_480)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2088_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i24_3_lut_4_lut_adj_328 (.A(bufcount[0]), .B(n30481), .C(rx_data[0]), 
         .D(\buffer[1] [0]), .Z(n11_adj_469)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_328.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_329 (.A(bufcount[0]), .B(n30481), .C(\buffer[1] [1]), 
         .D(rx_data[1]), .Z(n11_adj_470)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_329.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_330 (.A(bufcount[0]), .B(n30481), .C(rx_data[2]), 
         .D(\buffer[1] [2]), .Z(n11_adj_471)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_330.init = 16'hfd20;
    LUT4 i14578_4_lut (.A(\sendcount[3] ), .B(n9), .C(sendcount_c[2]), 
         .D(n30430), .Z(n3[3])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(271[10:37])
    defparam i14578_4_lut.init = 16'h4888;
    LUT4 i1_2_lut_3_lut_adj_331 (.A(n1295[3]), .B(n30375), .C(\buffer[2] [7]), 
         .Z(n28063)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_331.init = 16'h8080;
    LUT4 i1_3_lut_4_lut (.A(n1295[15]), .B(n9291), .C(n30383), .D(n1295[18]), 
         .Z(n13571)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_4_lut.init = 16'hf080;
    LUT4 i1_2_lut_3_lut_adj_332 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [0]), 
         .Z(n28071)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_332.init = 16'h8080;
    PFUMX i22358 (.BLUT(n30544), .ALUT(n30543), .C0(bufcount[2]), .Z(n30545));
    LUT4 i1_2_lut_3_lut_adj_333 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [1]), 
         .Z(n28069)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_333.init = 16'h8080;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n1295[15]), .B(n9291), .C(esc_data[1]), 
         .D(n1295[18]), .Z(n2037[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_3_lut_4_lut.init = 16'hf088;
    LUT4 i1_2_lut_3_lut_adj_334 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [2]), 
         .Z(n28070)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_334.init = 16'h8080;
    LUT4 i1_4_lut_adj_335 (.A(n5632), .B(n9297[0]), .C(n30383), .D(n1313), 
         .Z(n16120)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_335.init = 16'h8000;
    LUT4 i1_3_lut_4_lut_adj_336 (.A(n1295[15]), .B(n9291), .C(busy), .D(n1295[16]), 
         .Z(n10768)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_4_lut_adj_336.init = 16'h8f88;
    LUT4 i1_3_lut_3_lut_4_lut_adj_337 (.A(n1295[15]), .B(n9291), .C(esc_data[3]), 
         .D(n1295[18]), .Z(n22)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_3_lut_4_lut_adj_337.init = 16'hf088;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_476)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 i1_3_lut_3_lut_4_lut_adj_338 (.A(n1295[15]), .B(n9291), .C(esc_data[4]), 
         .D(n1295[18]), .Z(n2037[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_3_lut_4_lut_adj_338.init = 16'hf088;
    LUT4 i1_2_lut_3_lut_4_lut_adj_339 (.A(n1295[15]), .B(n9291), .C(n30383), 
         .D(n1295[18]), .Z(n18556)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_4_lut_adj_339.init = 16'h0080;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_474)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 i1_3_lut_3_lut_4_lut_adj_340 (.A(n1295[15]), .B(n9291), .C(esc_data[0]), 
         .D(n1295[18]), .Z(n2037[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_3_lut_4_lut_adj_340.init = 16'hf088;
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2621), .CK(debug_c_c), 
            .Q(register_addr_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_473)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2621), .CK(debug_c_c), 
            .Q(register_addr_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2621), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2621), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2621), .CK(debug_c_c), 
            .Q(register_addr[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2621), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2621), .CK(debug_c_c), 
            .Q(\register_addr[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_472)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 i9184_4_lut (.A(escape), .B(n12888), .C(n6_adj_481), .D(n1295[3]), 
         .Z(n10550)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i9184_4_lut.init = 16'h1aaa;
    LUT4 i2_2_lut_adj_341 (.A(debug_c_7), .B(n30383), .Z(n6_adj_481)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_341.init = 16'h8888;
    FD1P3IX buffer_0___i2 (.D(n27490), .SP(n9055), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_342 (.A(n27954), .B(rx_data[4]), .C(rx_data[1]), 
         .D(rx_data[3]), .Z(n12888)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i2_4_lut_adj_342.init = 16'hbfff;
    FD1P3IX buffer_0___i3 (.D(n27630), .SP(n9055), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n27494), .SP(n9055), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n27572), .SP(n9055), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n27506), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n27512), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n27508), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n27580), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n27576), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n27628), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n27504), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n27510), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n27574), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n27464), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n27586), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n26538), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n26541), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n26525), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n26535), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n26529), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i22 (.D(n26533), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    FD1P3IX buffer_0___i23 (.D(n26531), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n26534), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n26647), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n26523), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n26648), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n26502), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n26646), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n26560), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n26644), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n26673), .SP(n9055), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n26623), .SP(n14398), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n26583), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n26641), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n26639), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n26614), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n26637), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n26619), .SP(n14398), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n26622), .SP(n14398), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n26611), .SP(n14398), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n26640), .SP(n14398), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n26632), .SP(n14398), .CD(n30357), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n26576), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n26579), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n26593), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n26608), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n26600), .SP(n14398), .CD(n32388), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 equal_142_i13_2_lut (.A(rx_data[6]), .B(rx_data[7]), .Z(n13_adj_448)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(134[12:17])
    defparam equal_142_i13_2_lut.init = 16'heeee;
    FD1S3IX state_FSM_i2 (.D(n27778), .CK(debug_c_c), .CD(n32388), .Q(n1295[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n27666), .CK(debug_c_c), .CD(n32388), .Q(n1295[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n11905), .CK(debug_c_c), .CD(n30357), .Q(n1295[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n28005), .CK(debug_c_c), .CD(n32388), .Q(n1295[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n28232), .CK(debug_c_c), .CD(n32388), .Q(n1295[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1295[5]), .CK(debug_c_c), .CD(n32388), .Q(n1295[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1295[6]), .CK(debug_c_c), .CD(n32388), .Q(n1295[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1295[7]), .CK(debug_c_c), .CD(n32388), .Q(n1295[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1295[8]), .CK(debug_c_c), .CD(n32388), 
            .Q(n1295[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1400), .CK(debug_c_c), .CD(n32388), .Q(n1295[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1295[10]), .CK(debug_c_c), .CD(n32388), 
            .Q(n1295[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1295[11]), .CK(debug_c_c), .CD(n32388), 
            .Q(n1295[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1295[12]), .CK(debug_c_c), .CD(n32388), 
            .Q(n1295[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1406), .CK(debug_c_c), .CD(n32388), .Q(n1313));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1407), .CK(debug_c_c), .CD(n32388), .Q(n1295[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n10768), .CK(debug_c_c), .CD(n32388), .Q(n1295[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n11907), .CK(debug_c_c), .CD(n32388), .Q(n1310));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n26588), .CK(debug_c_c), .CD(n32388), .Q(n1295[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n10747), .CK(debug_c_c), .CD(n32388), .Q(n1295[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i21 (.D(n12021), .CK(debug_c_c), .CD(n32388), .Q(n1307));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5_rep_483 (.D(\buffer[1] [5]), .SP(n2621), .CK(debug_c_c), 
            .Q(n32377)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5_rep_483.GSR = "ENABLED";
    LUT4 i15257_3_lut_rep_350 (.A(n1295[13]), .B(n30383), .C(n1313), .Z(n30359)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15257_3_lut_rep_350.init = 16'hc8c8;
    LUT4 i21679_2_lut_3_lut (.A(n1295[13]), .B(n30383), .C(n1313), .Z(n9116)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i21679_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_adj_343 (.A(n1295[6]), .B(n1295[11]), .Z(n1748)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_343.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_344 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [3]), 
         .Z(n28060)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_344.init = 16'h8080;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n13571), .CD(n18556), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n13571), .CD(n18556), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_345 (.A(\buffer[0] [3]), .B(\buffer[0] [5]), .C(\buffer[0] [4]), 
         .D(\buffer[0] [6]), .Z(n12_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i3_4_lut_adj_345.init = 16'hfffe;
    LUT4 i21677_2_lut (.A(sendcount[0]), .B(n9), .Z(n21586)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i21677_2_lut.init = 16'h7777;
    LUT4 i1_2_lut_3_lut_adj_346 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [4]), 
         .Z(n28072)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_346.init = 16'h8080;
    LUT4 i1_4_lut_adj_347 (.A(sendcount_c[4]), .B(n5_adj_482), .C(n17), 
         .D(n4), .Z(n9)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_347.init = 16'hfffe;
    LUT4 i1_4_lut_adj_348 (.A(\reg_size[2] ), .B(sendcount_c[1]), .C(sendcount_c[2]), 
         .D(n30454), .Z(n5_adj_482)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C+(D))+!B !(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_348.init = 16'hed7b;
    LUT4 i1_4_lut_then_4_lut_adj_349 (.A(sendcount_c[4]), .B(sendcount[0]), 
         .C(sendcount_c[1]), .D(sendcount_c[2]), .Z(n30493)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut_adj_349.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_adj_350 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [5]), 
         .Z(n28074)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_350.init = 16'h8080;
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n13571), .CD(n18556), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n13571), .CD(n18556), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n13574), .CD(n16120), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n13574), .CD(n16120), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n13574), .CD(n16120), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n13574), .CD(n16120), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_351 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [6]), 
         .Z(n28073)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_351.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_352 (.A(n1295[3]), .B(n30375), .C(\buffer[3] [7]), 
         .Z(n28061)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_352.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_353 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [0]), 
         .Z(n28075)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_353.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_354 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [1]), 
         .Z(n28057)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_354.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_355 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [2]), 
         .Z(n28076)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_355.init = 16'h8080;
    LUT4 i1_2_lut_adj_356 (.A(\register_addr[1] ), .B(\steps_reg[7] ), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_356.init = 16'h8888;
    LUT4 i940_2_lut (.A(n1295[5]), .B(n30383), .Z(n2623)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i940_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_357 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [3]), 
         .Z(n28077)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_357.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_358 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [4]), 
         .Z(n28078)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_358.init = 16'h8080;
    LUT4 \buffer_0[[0__bdd_4_lut_22328  (.A(\buffer[0] [0]), .B(n28318), 
         .C(n15966), .D(n1748), .Z(n30297)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam \buffer_0[[0__bdd_4_lut_22328 .init = 16'h22f0;
    LUT4 \buffer_0[[0__bdd_4_lut  (.A(\buffer[0] [0]), .B(n28318), .C(n15968), 
         .D(n1748), .Z(n30298)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam \buffer_0[[0__bdd_4_lut .init = 16'h11f0;
    LUT4 i1_2_lut_3_lut_adj_359 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [5]), 
         .Z(n28079)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_359.init = 16'h8080;
    LUT4 i496_2_lut (.A(n1295[3]), .B(n1295[4]), .Z(n1696)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i496_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_360 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [6]), 
         .Z(n28080)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_360.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_361 (.A(n1295[3]), .B(n30375), .C(\buffer[4] [7]), 
         .Z(n28081)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_361.init = 16'h8080;
    LUT4 i1_4_lut_adj_362 (.A(esc_data[0]), .B(n30497), .C(esc_data[7]), 
         .D(esc_data[5]), .Z(n9291)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_362.init = 16'h0008;
    LUT4 i21436_4_lut (.A(rx_data[3]), .B(n30435), .C(rx_data[1]), .D(rx_data[4]), 
         .Z(n28589)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21436_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_363 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [0]), 
         .Z(n28082)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_363.init = 16'h8080;
    LUT4 i1_2_lut_adj_364 (.A(register_addr[0]), .B(\control_reg[7] ), .Z(n1_adj_216)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_364.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_365 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [1]), 
         .Z(n28083)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_365.init = 16'h8080;
    LUT4 i1_2_lut_adj_366 (.A(\register_addr[1] ), .B(\steps_reg[4] ), .Z(n17_adj_217)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_366.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_367 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [2]), 
         .Z(n28084)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_367.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_368 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [3]), 
         .Z(n28085)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_368.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_369 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [4]), 
         .Z(n28086)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_369.init = 16'h8080;
    LUT4 i14844_2_lut (.A(rx_data[2]), .B(rx_data[1]), .Z(n21219)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14844_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_370 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [5]), 
         .Z(n28088)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_370.init = 16'h8080;
    LUT4 i1_2_lut_adj_371 (.A(sendcount[0]), .B(\sendcount[3] ), .Z(n4_adj_218)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_371.init = 16'h4444;
    LUT4 i1_2_lut_adj_372 (.A(\register_addr[1] ), .B(\steps_reg[6] ), .Z(n13)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_372.init = 16'h8888;
    LUT4 i2_3_lut_rep_308_4_lut (.A(rw), .B(n30373), .C(n30417), .D(n28218), 
         .Z(n30317)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_308_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_adj_373 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [6]), 
         .Z(n28058)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_373.init = 16'h8080;
    LUT4 i1_2_lut_adj_374 (.A(\register_addr[1] ), .B(\steps_reg[5] ), .Z(n14)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_374.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_375 (.A(n1295[3]), .B(n30375), .C(\buffer[5] [7]), 
         .Z(n28087)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_375.init = 16'h8080;
    LUT4 i1_2_lut_adj_376 (.A(n1295[16]), .B(n1295[19]), .Z(n2046)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_376.init = 16'heeee;
    LUT4 i1_2_lut_adj_377 (.A(\register_addr[1] ), .B(\steps_reg[3] ), .Z(n12)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_377.init = 16'h8888;
    FD1P3AX rw_498_rep_485 (.D(n1295[10]), .SP(n2621), .CK(debug_c_c), 
            .Q(n32379));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_485.GSR = "ENABLED";
    LUT4 i21709_2_lut_2_lut (.A(n30383), .B(n9055), .Z(n14398)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21709_2_lut_2_lut.init = 16'hdddd;
    LUT4 i14459_2_lut (.A(\sendcount[3] ), .B(sendcount[0]), .Z(n9297[0])) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i14459_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_adj_378 (.A(register_addr[0]), .B(\control_reg[7]_adj_219 ), 
         .Z(n8263)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_378.init = 16'h4444;
    LUT4 i1_2_lut_adj_379 (.A(register_addr[0]), .B(\control_reg[7]_adj_220 ), 
         .Z(n8272)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_379.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_380 (.A(n1295[3]), .B(n30375), .C(n1295[13]), 
         .Z(n14_c)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_380.init = 16'hf8f8;
    PFUMX i22349 (.BLUT(n30522), .ALUT(n30523), .C0(sendcount[0]), .Z(n30524));
    PFUMX i22347 (.BLUT(n30519), .ALUT(n30520), .C0(sendcount[0]), .Z(n30521));
    PFUMX i22345 (.BLUT(n30516), .ALUT(n30517), .C0(sendcount[0]), .Z(n30518));
    PFUMX i22343 (.BLUT(n30513), .ALUT(n30514), .C0(sendcount[0]), .Z(n30515));
    LUT4 i1_2_lut_3_lut_adj_381 (.A(n1295[3]), .B(n30375), .C(\buffer[2] [0]), 
         .Z(n28064)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_381.init = 16'h8080;
    PFUMX i22341 (.BLUT(n30510), .ALUT(n30511), .C0(sendcount[0]), .Z(n30512));
    PFUMX i22339 (.BLUT(n30507), .ALUT(n30508), .C0(sendcount[0]), .Z(n30509));
    PFUMX i22337 (.BLUT(n30504), .ALUT(n30505), .C0(sendcount[0]), .Z(n30506));
    PFUMX i22335 (.BLUT(n30501), .ALUT(n30502), .C0(sendcount[0]), .Z(n30503));
    PFUMX i22333 (.BLUT(n30498), .ALUT(n30499), .C0(n30351), .Z(n30500));
    PFUMX i22331 (.BLUT(n30495), .ALUT(n30496), .C0(esc_data[2]), .Z(n30497));
    LUT4 i1_2_lut_3_lut_adj_382 (.A(n1295[3]), .B(n30375), .C(\buffer[2] [1]), 
         .Z(n28066)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_382.init = 16'h8080;
    PFUMX i22329 (.BLUT(n30492), .ALUT(n30493), .C0(\sendcount[3] ), .Z(n5632));
    \UARTTransmitter(baud_div=12)  uart_output (.n32388(n32388), .tx_data({tx_data}), 
            .send(send), .\reset_count[14] (\reset_count[14] ), .\reset_count[13] (\reset_count[13] ), 
            .\reset_count[12] (\reset_count[12] ), .n26787(n26787), .n30383(n30383), 
            .n30357(n30357), .busy(busy), .n10643(n10643), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_c(debug_c_c), .n30383(n30383), 
            .n32388(n32388), .n30357(n30357), .rx_data({rx_data}), .uart_rx_c(uart_rx_c), 
            .debug_c_7(debug_c_7), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (n32388, tx_data, send, \reset_count[14] , 
            \reset_count[13] , \reset_count[12] , n26787, n30383, n30357, 
            busy, n10643, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output n32388;
    input [7:0]tx_data;
    input send;
    input \reset_count[14] ;
    input \reset_count[13] ;
    input \reset_count[12] ;
    input n26787;
    output n30383;
    output n30357;
    output busy;
    output n10643;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n13441, n27434, n30204;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9037, n29553, n29554, n29545, n2, n17, n7, n10, n104, 
        n30202, n30203, n28257, n21151, n28607, n28608, n28609, 
        n30362, n2618, n28243, n28244, n2_adj_422;
    
    FD1P3AX state__i3 (.D(n27434), .SP(n13441), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n30204), .CK(bclk), .CD(n32388), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9037), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 n29553_bdd_2_lut (.A(n29553), .B(state[2]), .Z(n29554)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n29553_bdd_2_lut.init = 16'h2222;
    LUT4 n28091_bdd_4_lut (.A(state[3]), .B(state[1]), .C(send), .D(state[0]), 
         .Z(n29545)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam n28091_bdd_4_lut.init = 16'h7ffe;
    LUT4 i1_4_lut_rep_374 (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n26787), .Z(n30383)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i1_4_lut_rep_374.init = 16'heeea;
    LUT4 i53_1_lut_rep_348_4_lut (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n26787), .Z(n30357)) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i53_1_lut_rep_348_4_lut.init = 16'h1115;
    FD1P3IX busy_34 (.D(n2), .SP(n29554), .CD(n32388), .CK(bclk), .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    LUT4 state_2__bdd_2_lut (.A(state[0]), .B(state[3]), .Z(n30202)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_2__bdd_2_lut.init = 16'h1111;
    LUT4 state_2__bdd_4_lut_22497 (.A(state[0]), .B(state[3]), .C(state[1]), 
         .D(send), .Z(n30203)) /* synthesis lut_function=(A (B (C (D)))+!A (B+(C+(D)))) */ ;
    defparam state_2__bdd_4_lut_22497.init = 16'hd554;
    LUT4 state_2__bdd_4_lut_22272 (.A(send), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n29553)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)))) */ ;
    defparam state_2__bdd_4_lut_22272.init = 16'hc002;
    LUT4 i53_1_lut_rep_494 (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n26787), .Z(n32388)) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i53_1_lut_rep_494.init = 16'h1115;
    LUT4 i1_2_lut (.A(send), .B(state[3]), .Z(n28257)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i14776_2_lut (.A(state[1]), .B(state[0]), .Z(n21151)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14776_2_lut.init = 16'heeee;
    PFUMX i21456 (.BLUT(n28607), .ALUT(n28608), .C0(state[1]), .Z(n28609));
    LUT4 i1_3_lut_rep_353 (.A(n30383), .B(state[2]), .C(state[3]), .Z(n30362)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut_rep_353.init = 16'h2a2a;
    LUT4 i1_3_lut_4_lut (.A(n30383), .B(state[2]), .C(state[3]), .D(n2618), 
         .Z(n28243)) /* synthesis lut_function=(!((B (C+(D))+!B !(D))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2208;
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9037), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9037), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9037), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9037), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9037), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9037), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9037), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    PFUMX i22273 (.BLUT(n30203), .ALUT(n30202), .C0(state[2]), .Z(n30204));
    LUT4 i1_3_lut (.A(state[1]), .B(n30362), .C(state[0]), .Z(n28244)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    LUT4 status_led_c_bdd_2_lut_22058_3_lut (.A(n30383), .B(state[2]), .C(n29545), 
         .Z(n13441)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam status_led_c_bdd_2_lut_22058_3_lut.init = 16'hfdfd;
    LUT4 i2_3_lut_4_lut (.A(n30383), .B(state[2]), .C(n21151), .D(n28257), 
         .Z(n9037)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0200;
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n32388), .CK(bclk), .Q(n10643)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i3_1_lut (.A(state[3]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i3_1_lut.init = 16'h5555;
    LUT4 i1_4_lut (.A(n30383), .B(state[3]), .C(state[2]), .D(n2618), 
         .Z(n27434)) /* synthesis lut_function=(!((B (C)+!B !(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h2808;
    LUT4 Mux_22_i7_4_lut (.A(n2_adj_422), .B(n28609), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2_adj_422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i14896_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i14896_4_lut.init = 16'hfcee;
    FD1P3AX state__i1 (.D(n28244), .SP(n13441), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX state__i2 (.D(n28243), .SP(n13441), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    LUT4 i935_2_lut (.A(state[0]), .B(state[1]), .Z(n2618)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i935_2_lut.init = 16'h8888;
    LUT4 i21454_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n28607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21454_3_lut.init = 16'hcaca;
    LUT4 i21455_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n28608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21455_3_lut.init = 16'hcaca;
    \ClockDividerP(factor=12)  baud_gen (.debug_c_c(debug_c_c), .GND_net(GND_net), 
            .bclk(bclk)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (debug_c_c, GND_net, bclk) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input GND_net;
    output bclk;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n16172;
    wire [31:0]n102;
    
    wire n26166, n8094, n26165, n26164, n26163, n26162, n26161, 
        n26160, n26159, n26158, n26157, n26156, n26155, n26154, 
        n26153, n26152, n26151, n28789, n49, n56, n50, n54, 
        n46, n28455, n52, n42, n48, n34, n26118, n26117, n26116, 
        n26115, n26114, n26113, n26112, n26111, n26110, n26109, 
        n26108, n26107, n26106, n26105, n26104, n26103;
    
    FD1S3IX count_2616__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i0.GSR = "ENABLED";
    CCU2D sub_2036_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26166), .S0(n8094));
    defparam sub_2036_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2036_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2036_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2036_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26165), .COUT(n26166));
    defparam sub_2036_add_2_32.INIT0 = 16'h5555;
    defparam sub_2036_add_2_32.INIT1 = 16'h5555;
    defparam sub_2036_add_2_32.INJECT1_0 = "NO";
    defparam sub_2036_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26164), .COUT(n26165));
    defparam sub_2036_add_2_30.INIT0 = 16'h5555;
    defparam sub_2036_add_2_30.INIT1 = 16'h5555;
    defparam sub_2036_add_2_30.INJECT1_0 = "NO";
    defparam sub_2036_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26163), .COUT(n26164));
    defparam sub_2036_add_2_28.INIT0 = 16'h5555;
    defparam sub_2036_add_2_28.INIT1 = 16'h5555;
    defparam sub_2036_add_2_28.INJECT1_0 = "NO";
    defparam sub_2036_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26162), .COUT(n26163));
    defparam sub_2036_add_2_26.INIT0 = 16'h5555;
    defparam sub_2036_add_2_26.INIT1 = 16'h5555;
    defparam sub_2036_add_2_26.INJECT1_0 = "NO";
    defparam sub_2036_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26161), .COUT(n26162));
    defparam sub_2036_add_2_24.INIT0 = 16'h5555;
    defparam sub_2036_add_2_24.INIT1 = 16'h5555;
    defparam sub_2036_add_2_24.INJECT1_0 = "NO";
    defparam sub_2036_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26160), .COUT(n26161));
    defparam sub_2036_add_2_22.INIT0 = 16'h5555;
    defparam sub_2036_add_2_22.INIT1 = 16'h5555;
    defparam sub_2036_add_2_22.INJECT1_0 = "NO";
    defparam sub_2036_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26159), .COUT(n26160));
    defparam sub_2036_add_2_20.INIT0 = 16'h5555;
    defparam sub_2036_add_2_20.INIT1 = 16'h5555;
    defparam sub_2036_add_2_20.INJECT1_0 = "NO";
    defparam sub_2036_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26158), .COUT(n26159));
    defparam sub_2036_add_2_18.INIT0 = 16'h5555;
    defparam sub_2036_add_2_18.INIT1 = 16'h5555;
    defparam sub_2036_add_2_18.INJECT1_0 = "NO";
    defparam sub_2036_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26157), .COUT(n26158));
    defparam sub_2036_add_2_16.INIT0 = 16'h5555;
    defparam sub_2036_add_2_16.INIT1 = 16'h5555;
    defparam sub_2036_add_2_16.INJECT1_0 = "NO";
    defparam sub_2036_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26156), .COUT(n26157));
    defparam sub_2036_add_2_14.INIT0 = 16'h5555;
    defparam sub_2036_add_2_14.INIT1 = 16'h5555;
    defparam sub_2036_add_2_14.INJECT1_0 = "NO";
    defparam sub_2036_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26155), .COUT(n26156));
    defparam sub_2036_add_2_12.INIT0 = 16'h5555;
    defparam sub_2036_add_2_12.INIT1 = 16'h5555;
    defparam sub_2036_add_2_12.INJECT1_0 = "NO";
    defparam sub_2036_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26154), .COUT(n26155));
    defparam sub_2036_add_2_10.INIT0 = 16'h5555;
    defparam sub_2036_add_2_10.INIT1 = 16'h5555;
    defparam sub_2036_add_2_10.INJECT1_0 = "NO";
    defparam sub_2036_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26153), .COUT(n26154));
    defparam sub_2036_add_2_8.INIT0 = 16'h5555;
    defparam sub_2036_add_2_8.INIT1 = 16'h5555;
    defparam sub_2036_add_2_8.INJECT1_0 = "NO";
    defparam sub_2036_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26152), .COUT(n26153));
    defparam sub_2036_add_2_6.INIT0 = 16'h5555;
    defparam sub_2036_add_2_6.INIT1 = 16'h5555;
    defparam sub_2036_add_2_6.INJECT1_0 = "NO";
    defparam sub_2036_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26151), .COUT(n26152));
    defparam sub_2036_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2036_add_2_4.INIT1 = 16'h5555;
    defparam sub_2036_add_2_4.INJECT1_0 = "NO";
    defparam sub_2036_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26151));
    defparam sub_2036_add_2_2.INIT0 = 16'h0000;
    defparam sub_2036_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2036_add_2_2.INJECT1_0 = "NO";
    defparam sub_2036_add_2_2.INJECT1_1 = "NO";
    FD1S3AX clk_o_14 (.D(n8094), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    LUT4 i21739_4_lut (.A(n28789), .B(n49), .C(n56), .D(n50), .Z(n16172)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21739_4_lut.init = 16'h0002;
    LUT4 i21737_4_lut (.A(count[31]), .B(n54), .C(n46), .D(n28455), 
         .Z(n28789)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21737_4_lut.init = 16'h0100;
    LUT4 i19_4_lut (.A(count[24]), .B(count[27]), .C(count[4]), .D(count[30]), 
         .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(count[5]), .B(n52), .C(n42), .D(count[6]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i20_4_lut (.A(count[7]), .B(count[19]), .C(count[14]), .D(count[22]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(count[16]), .B(n48), .C(n34), .D(count[11]), 
         .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(count[28]), .B(count[2]), .C(count[18]), .D(count[8]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i21308_3_lut (.A(count[3]), .B(count[0]), .C(count[1]), .Z(n28455)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i21308_3_lut.init = 16'h8080;
    LUT4 i18_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[21]), .B(count[25]), .Z(n34)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(count[15]), .B(count[29]), .C(count[23]), .D(count[13]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i12_2_lut (.A(count[10]), .B(count[20]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i12_2_lut.init = 16'heeee;
    CCU2D count_2616_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26118), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_33.INIT1 = 16'h0000;
    defparam count_2616_add_4_33.INJECT1_0 = "NO";
    defparam count_2616_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26117), .COUT(n26118), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_31.INJECT1_0 = "NO";
    defparam count_2616_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26116), .COUT(n26117), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_29.INJECT1_0 = "NO";
    defparam count_2616_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26115), .COUT(n26116), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_27.INJECT1_0 = "NO";
    defparam count_2616_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26114), .COUT(n26115), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_25.INJECT1_0 = "NO";
    defparam count_2616_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26113), .COUT(n26114), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_23.INJECT1_0 = "NO";
    defparam count_2616_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26112), .COUT(n26113), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_21.INJECT1_0 = "NO";
    defparam count_2616_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26111), .COUT(n26112), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_19.INJECT1_0 = "NO";
    defparam count_2616_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26110), .COUT(n26111), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_17.INJECT1_0 = "NO";
    defparam count_2616_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26109), .COUT(n26110), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_15.INJECT1_0 = "NO";
    defparam count_2616_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26108), .COUT(n26109), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_13.INJECT1_0 = "NO";
    defparam count_2616_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26107), .COUT(n26108), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_11.INJECT1_0 = "NO";
    defparam count_2616_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26106), .COUT(n26107), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_9.INJECT1_0 = "NO";
    defparam count_2616_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26105), .COUT(n26106), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_7.INJECT1_0 = "NO";
    defparam count_2616_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26104), .COUT(n26105), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_5.INJECT1_0 = "NO";
    defparam count_2616_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26103), .COUT(n26104), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2616_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2616_add_4_3.INJECT1_0 = "NO";
    defparam count_2616_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2616_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26103), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616_add_4_1.INIT0 = 16'hF000;
    defparam count_2616_add_4_1.INIT1 = 16'h0555;
    defparam count_2616_add_4_1.INJECT1_0 = "NO";
    defparam count_2616_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2616__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i1.GSR = "ENABLED";
    FD1S3IX count_2616__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i2.GSR = "ENABLED";
    FD1S3IX count_2616__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i3.GSR = "ENABLED";
    FD1S3IX count_2616__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i4.GSR = "ENABLED";
    FD1S3IX count_2616__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i5.GSR = "ENABLED";
    FD1S3IX count_2616__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i6.GSR = "ENABLED";
    FD1S3IX count_2616__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i7.GSR = "ENABLED";
    FD1S3IX count_2616__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i8.GSR = "ENABLED";
    FD1S3IX count_2616__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i9.GSR = "ENABLED";
    FD1S3IX count_2616__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i10.GSR = "ENABLED";
    FD1S3IX count_2616__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i11.GSR = "ENABLED";
    FD1S3IX count_2616__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i12.GSR = "ENABLED";
    FD1S3IX count_2616__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i13.GSR = "ENABLED";
    FD1S3IX count_2616__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i14.GSR = "ENABLED";
    FD1S3IX count_2616__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i15.GSR = "ENABLED";
    FD1S3IX count_2616__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i16.GSR = "ENABLED";
    FD1S3IX count_2616__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i17.GSR = "ENABLED";
    FD1S3IX count_2616__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i18.GSR = "ENABLED";
    FD1S3IX count_2616__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i19.GSR = "ENABLED";
    FD1S3IX count_2616__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i20.GSR = "ENABLED";
    FD1S3IX count_2616__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i21.GSR = "ENABLED";
    FD1S3IX count_2616__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i22.GSR = "ENABLED";
    FD1S3IX count_2616__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i23.GSR = "ENABLED";
    FD1S3IX count_2616__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i24.GSR = "ENABLED";
    FD1S3IX count_2616__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i25.GSR = "ENABLED";
    FD1S3IX count_2616__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i26.GSR = "ENABLED";
    FD1S3IX count_2616__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i27.GSR = "ENABLED";
    FD1S3IX count_2616__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i28.GSR = "ENABLED";
    FD1S3IX count_2616__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i29.GSR = "ENABLED";
    FD1S3IX count_2616__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i30.GSR = "ENABLED";
    FD1S3IX count_2616__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16172), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2616__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_c, n30383, n32388, n30357, 
            rx_data, uart_rx_c, debug_c_7, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30383;
    input n32388;
    input n30357;
    output [7:0]rx_data;
    input uart_rx_c;
    output debug_c_7;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n32;
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n30424, bclk, n27460;
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n9013, n27066, n29536, n15173, n27388, n32374, n9027, 
        n9025, n9023, n9021, n9019, n9017, n9015, n9011, n9009, 
        n9007, n9005, n9003, n9001, n8985, n8987, baud_reset, 
        n19;
    wire [7:0]n78;
    
    wire n13059, n13, n28294, n30462, n28352, n25, n27, n30441, 
        n30451, n30409, n30836, n30835, n29, n15172, n21, n23, 
        n28550, n21_adj_417, n30410, n29535, n30464, n30452, n28334, 
        n25_adj_418, n19_adj_419, n21519, n30465, n13068, n19_adj_420, 
        n4, n29534, n33;
    wire [5:0]n6;
    
    wire n4_adj_421;
    
    LUT4 i1_2_lut_rep_415 (.A(n32), .B(state[5]), .Z(n30424)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_415.init = 16'h2222;
    LUT4 i1_3_lut_4_lut (.A(n32), .B(state[5]), .C(state[0]), .D(bclk), 
         .Z(n27460)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut.init = 16'hf200;
    FD1P3AX rdata_i0_i7 (.D(n9013), .SP(n30383), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n27066), .CK(debug_c_c), .CD(n32388), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n29536), .CK(debug_c_c), .CD(n32388), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n15173), .CK(debug_c_c), .CD(n30357), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n27388), .CK(debug_c_c), .CD(n30357), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n32374), .CK(debug_c_c), .CD(n30357), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n9027), .SP(n30383), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n9025), .SP(n30383), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n9023), .SP(n30383), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n9021), .SP(n30383), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n9019), .SP(n30383), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n9017), .SP(n30383), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n9015), .SP(n30383), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n9011), .SP(n30383), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n9009), .SP(n30383), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n9007), .SP(n30383), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n9005), .SP(n30383), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n9003), .SP(n30383), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i1 (.D(n9001), .SP(n30383), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i0 (.D(n8985), .SP(n30383), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n8987), .SP(n30383), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n27460), .CK(debug_c_c), .CD(n30357), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n19), .CK(debug_c_c), .PD(n32388), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n78[4]), .B(rdata[4]), .C(n13059), .D(n13), .Z(n9007)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i4327_4_lut (.A(uart_rx_c), .B(rdata[4]), .C(state[2]), .D(n28294), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4327_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_210 (.A(n78[3]), .B(rdata[3]), .C(n13059), .D(n13), 
         .Z(n9005)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_210.init = 16'heca0;
    LUT4 i4332_4_lut (.A(uart_rx_c), .B(rdata[3]), .C(n30462), .D(n28352), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4332_4_lut.init = 16'hccac;
    LUT4 i1_2_lut (.A(state[3]), .B(state[2]), .Z(n28352)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut.init = 16'hbbbb;
    PFUMX i40 (.BLUT(n25), .ALUT(n27), .C0(state[0]), .Z(n27388));
    LUT4 i1_4_lut_adj_211 (.A(n78[2]), .B(rdata[2]), .C(n13059), .D(n13), 
         .Z(n9003)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_211.init = 16'heca0;
    LUT4 i4334_4_lut (.A(uart_rx_c), .B(rdata[2]), .C(n30441), .D(n28352), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4334_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_212 (.A(n78[1]), .B(rdata[1]), .C(n13059), .D(n13), 
         .Z(n9001)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_212.init = 16'heca0;
    LUT4 i4336_4_lut (.A(uart_rx_c), .B(rdata[1]), .C(n30451), .D(n30462), 
         .Z(n78[1])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4336_4_lut.init = 16'hcacc;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(n30409), .C(n32), .D(uart_rx_c), 
         .Z(n30836)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+(D))) */ ;
    defparam state_1__bdd_4_lut.init = 16'ha2b3;
    LUT4 state_1__bdd_2_lut (.A(state[1]), .B(bclk), .Z(n30835)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam state_1__bdd_2_lut.init = 16'h9999;
    PFUMX i8761 (.BLUT(n29), .ALUT(n15172), .C0(state[0]), .Z(n15173));
    PFUMX i36 (.BLUT(n21), .ALUT(n23), .C0(state[5]), .Z(n27066));
    LUT4 n30836_bdd_4_lut (.A(n30836), .B(state[5]), .C(n30835), .D(state[0]), 
         .Z(n32374)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam n30836_bdd_4_lut.init = 16'hf022;
    LUT4 i1_4_lut_adj_213 (.A(state[5]), .B(n28550), .C(state[2]), .D(n21_adj_417), 
         .Z(n25)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_213.init = 16'h5111;
    LUT4 i1_2_lut_rep_432 (.A(state[1]), .B(bclk), .Z(n30441)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_rep_432.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut (.A(state[1]), .B(bclk), .C(state[3]), .Z(n28294)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i41_3_lut (.A(state[1]), .B(state[2]), .C(bclk), .Z(n27)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i41_3_lut.init = 16'hc6c6;
    LUT4 n28089_bdd_4_lut (.A(n30424), .B(state[4]), .C(bclk), .D(n30410), 
         .Z(n29535)) /* synthesis lut_function=(!((B (C (D))+!B !(C (D)))+!A)) */ ;
    defparam n28089_bdd_4_lut.init = 16'h2888;
    LUT4 i2_2_lut_rep_442 (.A(state[3]), .B(state[2]), .Z(n30451)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_2_lut_rep_442.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[3]), .B(state[2]), .C(n30464), 
         .D(n30452), .Z(n28334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_214 (.A(state[3]), .B(state[2]), .C(n30452), 
         .D(state[0]), .Z(n25_adj_418)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut_adj_214.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_215 (.A(state[3]), .B(state[2]), .C(n32), 
         .D(n30452), .Z(n21_adj_417)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut_adj_215.init = 16'hf0f1;
    LUT4 i21397_2_lut_3_lut_4_lut (.A(state[3]), .B(state[2]), .C(uart_rx_c), 
         .D(n30452), .Z(n28550)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21397_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_443 (.A(state[1]), .B(state[4]), .Z(n30452)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_443.init = 16'heeee;
    LUT4 i2_2_lut_rep_400_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(state[2]), 
         .D(state[3]), .Z(n30409)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_2_lut_rep_400_3_lut_4_lut.init = 16'hfffe;
    FD1S3IX drdy_51 (.D(n19_adj_419), .CK(debug_c_c), .CD(n32388), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 i14523_2_lut_rep_453 (.A(bclk), .B(state[1]), .Z(n30462)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14523_2_lut_rep_453.init = 16'h8888;
    LUT4 i15141_2_lut_3_lut (.A(bclk), .B(state[1]), .C(state[3]), .Z(n21519)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15141_2_lut_3_lut.init = 16'h8080;
    LUT4 i14416_2_lut_rep_455 (.A(state[0]), .B(state[5]), .Z(n30464)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14416_2_lut_rep_455.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_216 (.A(state[0]), .B(state[5]), .C(state[4]), 
         .Z(n13059)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_216.init = 16'h1010;
    LUT4 i3374_3_lut_rep_456 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n30465)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3374_3_lut_rep_456.init = 16'h8080;
    LUT4 i3381_2_lut_rep_401_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n30410)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3381_2_lut_rep_401_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_217 (.A(n78[0]), .B(rdata[0]), .C(n13059), .D(n13), 
         .Z(n8985)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_217.init = 16'heca0;
    LUT4 i4370_4_lut (.A(uart_rx_c), .B(rdata[0]), .C(n30451), .D(n30441), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4370_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_218 (.A(rdata[0]), .B(rx_data[0]), .C(n13068), .D(n19_adj_420), 
         .Z(n8987)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_218.init = 16'heca0;
    LUT4 i1_4_lut_adj_219 (.A(state[4]), .B(state[3]), .C(state[2]), .D(state[1]), 
         .Z(n32)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_219.init = 16'heaaa;
    LUT4 i2_3_lut_4_lut (.A(n30452), .B(n30451), .C(state[0]), .D(state[5]), 
         .Z(n13068)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_4_lut_adj_220 (.A(n30452), .B(n30451), .C(state[0]), 
         .D(state[5]), .Z(n19_adj_420)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i2_3_lut_4_lut_adj_220.init = 16'hfeff;
    LUT4 i21747_4_lut (.A(baud_reset), .B(n28334), .C(uart_rx_c), .D(n25_adj_418), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21747_4_lut.init = 16'ha8ec;
    LUT4 i1_2_lut_3_lut_adj_221 (.A(state[3]), .B(n30465), .C(state[4]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_221.init = 16'h8080;
    LUT4 n28089_bdd_3_lut_4_lut (.A(state[3]), .B(n30465), .C(bclk), .D(state[4]), 
         .Z(n29534)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n28089_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 i1_4_lut_4_lut (.A(state[3]), .B(n30465), .C(bclk), .D(n32), 
         .Z(n33)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h6a00;
    LUT4 i8760_3_lut_3_lut (.A(state[3]), .B(n30465), .C(bclk), .Z(n15172)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i8760_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i1_4_lut_adj_222 (.A(n78[6]), .B(rdata[6]), .C(n13059), .D(n13), 
         .Z(n9011)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_222.init = 16'heca0;
    LUT4 i4323_4_lut (.A(uart_rx_c), .B(rdata[6]), .C(state[2]), .D(n28294), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4323_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_223 (.A(n78[7]), .B(rdata[7]), .C(n13059), .D(n13), 
         .Z(n9013)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_223.init = 16'heca0;
    LUT4 i4321_4_lut (.A(rdata[7]), .B(uart_rx_c), .C(state[2]), .D(n21519), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4321_4_lut.init = 16'hcaaa;
    LUT4 i21326_4_lut (.A(n6[3]), .B(state[5]), .C(n33), .D(n30409), 
         .Z(n29)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21326_4_lut.init = 16'h3032;
    LUT4 i14462_2_lut (.A(state[3]), .B(uart_rx_c), .Z(n6[3])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(42[8] 47[12])
    defparam i14462_2_lut.init = 16'hbbbb;
    LUT4 i2_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut.init = 16'hefef;
    LUT4 i2_4_lut (.A(bclk), .B(n4), .C(state[0]), .D(n32), .Z(n21)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'h4840;
    LUT4 i38_4_lut (.A(n28550), .B(n30410), .C(state[0]), .D(n4_adj_421), 
         .Z(n23)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i38_4_lut.init = 16'hf535;
    LUT4 i1_2_lut_adj_224 (.A(state[4]), .B(bclk), .Z(n4_adj_421)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_224.init = 16'hdddd;
    LUT4 i1_4_lut_adj_225 (.A(n78[5]), .B(rdata[5]), .C(n13059), .D(n13), 
         .Z(n9009)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_225.init = 16'heca0;
    LUT4 i4325_4_lut (.A(uart_rx_c), .B(rdata[5]), .C(state[2]), .D(n21519), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4325_4_lut.init = 16'hcacc;
    PFUMX i22014 (.BLUT(n29535), .ALUT(n29534), .C0(state[0]), .Z(n29536));
    LUT4 i1_4_lut_adj_226 (.A(rdata[7]), .B(rx_data[7]), .C(n13068), .D(n19_adj_420), 
         .Z(n9027)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_226.init = 16'heca0;
    LUT4 i21745_4_lut (.A(debug_c_7), .B(n28334), .C(uart_rx_c), .D(n25_adj_418), 
         .Z(n19_adj_419)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21745_4_lut.init = 16'ha8ec;
    LUT4 i1_4_lut_adj_227 (.A(rdata[6]), .B(rx_data[6]), .C(n13068), .D(n19_adj_420), 
         .Z(n9025)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_227.init = 16'heca0;
    LUT4 i1_4_lut_adj_228 (.A(rdata[5]), .B(rx_data[5]), .C(n13068), .D(n19_adj_420), 
         .Z(n9023)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_228.init = 16'heca0;
    LUT4 i1_4_lut_adj_229 (.A(rdata[4]), .B(rx_data[4]), .C(n13068), .D(n19_adj_420), 
         .Z(n9021)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_229.init = 16'heca0;
    LUT4 i1_4_lut_adj_230 (.A(rdata[3]), .B(rx_data[3]), .C(n13068), .D(n19_adj_420), 
         .Z(n9019)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_230.init = 16'heca0;
    LUT4 i1_4_lut_adj_231 (.A(rdata[2]), .B(rx_data[2]), .C(n13068), .D(n19_adj_420), 
         .Z(n9017)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_231.init = 16'heca0;
    LUT4 i1_4_lut_adj_232 (.A(rdata[1]), .B(rx_data[1]), .C(n13068), .D(n19_adj_420), 
         .Z(n9015)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_232.init = 16'heca0;
    \ClockDividerP(factor=12)_U0  baud_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .bclk(bclk), .baud_reset(baud_reset)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (GND_net, debug_c_c, bclk, baud_reset) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    output bclk;
    input baud_reset;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n26198, n8059, n26197;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n26196, n26195, n26194, n26193, n26192, n26191, n26190, 
        n26189, n26188, n26187, n26186, n26185, n26184, n26183, 
        n2773;
    wire [31:0]n134;
    
    wire n26102, n26101, n26100, n26099, n26098, n26097, n26096, 
        n26095, n26094, n26093, n26092, n26091, n26090, n26089, 
        n26088, n26087, n55, n26392, n56, n52, n44, n35, n54, 
        n48, n36, n46, n32, n50, n40;
    
    CCU2D sub_2034_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26198), .S0(n8059));
    defparam sub_2034_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2034_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2034_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2034_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26197), .COUT(n26198));
    defparam sub_2034_add_2_32.INIT0 = 16'h5555;
    defparam sub_2034_add_2_32.INIT1 = 16'h5555;
    defparam sub_2034_add_2_32.INJECT1_0 = "NO";
    defparam sub_2034_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26196), .COUT(n26197));
    defparam sub_2034_add_2_30.INIT0 = 16'h5555;
    defparam sub_2034_add_2_30.INIT1 = 16'h5555;
    defparam sub_2034_add_2_30.INJECT1_0 = "NO";
    defparam sub_2034_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26195), .COUT(n26196));
    defparam sub_2034_add_2_28.INIT0 = 16'h5555;
    defparam sub_2034_add_2_28.INIT1 = 16'h5555;
    defparam sub_2034_add_2_28.INJECT1_0 = "NO";
    defparam sub_2034_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26194), .COUT(n26195));
    defparam sub_2034_add_2_26.INIT0 = 16'h5555;
    defparam sub_2034_add_2_26.INIT1 = 16'h5555;
    defparam sub_2034_add_2_26.INJECT1_0 = "NO";
    defparam sub_2034_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26193), .COUT(n26194));
    defparam sub_2034_add_2_24.INIT0 = 16'h5555;
    defparam sub_2034_add_2_24.INIT1 = 16'h5555;
    defparam sub_2034_add_2_24.INJECT1_0 = "NO";
    defparam sub_2034_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26192), .COUT(n26193));
    defparam sub_2034_add_2_22.INIT0 = 16'h5555;
    defparam sub_2034_add_2_22.INIT1 = 16'h5555;
    defparam sub_2034_add_2_22.INJECT1_0 = "NO";
    defparam sub_2034_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26191), .COUT(n26192));
    defparam sub_2034_add_2_20.INIT0 = 16'h5555;
    defparam sub_2034_add_2_20.INIT1 = 16'h5555;
    defparam sub_2034_add_2_20.INJECT1_0 = "NO";
    defparam sub_2034_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26190), .COUT(n26191));
    defparam sub_2034_add_2_18.INIT0 = 16'h5555;
    defparam sub_2034_add_2_18.INIT1 = 16'h5555;
    defparam sub_2034_add_2_18.INJECT1_0 = "NO";
    defparam sub_2034_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26189), .COUT(n26190));
    defparam sub_2034_add_2_16.INIT0 = 16'h5555;
    defparam sub_2034_add_2_16.INIT1 = 16'h5555;
    defparam sub_2034_add_2_16.INJECT1_0 = "NO";
    defparam sub_2034_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26188), .COUT(n26189));
    defparam sub_2034_add_2_14.INIT0 = 16'h5555;
    defparam sub_2034_add_2_14.INIT1 = 16'h5555;
    defparam sub_2034_add_2_14.INJECT1_0 = "NO";
    defparam sub_2034_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26187), .COUT(n26188));
    defparam sub_2034_add_2_12.INIT0 = 16'h5555;
    defparam sub_2034_add_2_12.INIT1 = 16'h5555;
    defparam sub_2034_add_2_12.INJECT1_0 = "NO";
    defparam sub_2034_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26186), .COUT(n26187));
    defparam sub_2034_add_2_10.INIT0 = 16'h5555;
    defparam sub_2034_add_2_10.INIT1 = 16'h5555;
    defparam sub_2034_add_2_10.INJECT1_0 = "NO";
    defparam sub_2034_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26185), .COUT(n26186));
    defparam sub_2034_add_2_8.INIT0 = 16'h5555;
    defparam sub_2034_add_2_8.INIT1 = 16'h5555;
    defparam sub_2034_add_2_8.INJECT1_0 = "NO";
    defparam sub_2034_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26184), .COUT(n26185));
    defparam sub_2034_add_2_6.INIT0 = 16'h5555;
    defparam sub_2034_add_2_6.INIT1 = 16'h5555;
    defparam sub_2034_add_2_6.INJECT1_0 = "NO";
    defparam sub_2034_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26183), .COUT(n26184));
    defparam sub_2034_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2034_add_2_4.INIT1 = 16'h5555;
    defparam sub_2034_add_2_4.INJECT1_0 = "NO";
    defparam sub_2034_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26183));
    defparam sub_2034_add_2_2.INIT0 = 16'h0000;
    defparam sub_2034_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2034_add_2_2.INJECT1_0 = "NO";
    defparam sub_2034_add_2_2.INJECT1_1 = "NO";
    FD1S3IX count_2615__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2773), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i0.GSR = "ENABLED";
    FD1S3IX clk_o_14 (.D(n8059), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2615_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26102), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_33.INIT1 = 16'h0000;
    defparam count_2615_add_4_33.INJECT1_0 = "NO";
    defparam count_2615_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26101), .COUT(n26102), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_31.INJECT1_0 = "NO";
    defparam count_2615_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26100), .COUT(n26101), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_29.INJECT1_0 = "NO";
    defparam count_2615_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26099), .COUT(n26100), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_27.INJECT1_0 = "NO";
    defparam count_2615_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26098), .COUT(n26099), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_25.INJECT1_0 = "NO";
    defparam count_2615_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26097), .COUT(n26098), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_23.INJECT1_0 = "NO";
    defparam count_2615_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26096), .COUT(n26097), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_21.INJECT1_0 = "NO";
    defparam count_2615_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26095), .COUT(n26096), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_19.INJECT1_0 = "NO";
    defparam count_2615_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26094), .COUT(n26095), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_17.INJECT1_0 = "NO";
    defparam count_2615_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26093), .COUT(n26094), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_15.INJECT1_0 = "NO";
    defparam count_2615_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26092), .COUT(n26093), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_13.INJECT1_0 = "NO";
    defparam count_2615_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26091), .COUT(n26092), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_11.INJECT1_0 = "NO";
    defparam count_2615_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26090), .COUT(n26091), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_9.INJECT1_0 = "NO";
    defparam count_2615_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26089), .COUT(n26090), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_7.INJECT1_0 = "NO";
    defparam count_2615_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26088), .COUT(n26089), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_5.INJECT1_0 = "NO";
    defparam count_2615_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26087), .COUT(n26088), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2615_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2615_add_4_3.INJECT1_0 = "NO";
    defparam count_2615_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2615_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26087), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615_add_4_1.INIT0 = 16'hF000;
    defparam count_2615_add_4_1.INIT1 = 16'h0555;
    defparam count_2615_add_4_1.INJECT1_0 = "NO";
    defparam count_2615_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2615__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2773), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i1.GSR = "ENABLED";
    FD1S3IX count_2615__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2773), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i2.GSR = "ENABLED";
    FD1S3IX count_2615__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2773), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i3.GSR = "ENABLED";
    FD1S3IX count_2615__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2773), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i4.GSR = "ENABLED";
    FD1S3IX count_2615__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2773), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i5.GSR = "ENABLED";
    FD1S3IX count_2615__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2773), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i6.GSR = "ENABLED";
    FD1S3IX count_2615__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2773), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i7.GSR = "ENABLED";
    FD1S3IX count_2615__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2773), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i8.GSR = "ENABLED";
    FD1S3IX count_2615__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2773), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i9.GSR = "ENABLED";
    FD1S3IX count_2615__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i10.GSR = "ENABLED";
    FD1S3IX count_2615__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i11.GSR = "ENABLED";
    FD1S3IX count_2615__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i12.GSR = "ENABLED";
    FD1S3IX count_2615__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i13.GSR = "ENABLED";
    FD1S3IX count_2615__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i14.GSR = "ENABLED";
    FD1S3IX count_2615__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i15.GSR = "ENABLED";
    FD1S3IX count_2615__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i16.GSR = "ENABLED";
    FD1S3IX count_2615__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i17.GSR = "ENABLED";
    FD1S3IX count_2615__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i18.GSR = "ENABLED";
    FD1S3IX count_2615__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i19.GSR = "ENABLED";
    FD1S3IX count_2615__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i20.GSR = "ENABLED";
    FD1S3IX count_2615__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i21.GSR = "ENABLED";
    FD1S3IX count_2615__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i22.GSR = "ENABLED";
    FD1S3IX count_2615__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i23.GSR = "ENABLED";
    FD1S3IX count_2615__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i24.GSR = "ENABLED";
    FD1S3IX count_2615__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i25.GSR = "ENABLED";
    FD1S3IX count_2615__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i26.GSR = "ENABLED";
    FD1S3IX count_2615__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i27.GSR = "ENABLED";
    FD1S3IX count_2615__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i28.GSR = "ENABLED";
    FD1S3IX count_2615__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i29.GSR = "ENABLED";
    FD1S3IX count_2615__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i30.GSR = "ENABLED";
    FD1S3IX count_2615__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2773), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2615__i31.GSR = "ENABLED";
    LUT4 i1090_4_lut (.A(n55), .B(baud_reset), .C(n26392), .D(n56), 
         .Z(n2773)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i1090_4_lut.init = 16'hccdc;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(count[1]), .B(count[3]), .C(count[0]), .Z(n26392)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (debug_c_c, n8894, n32384, 
            databus, n608, n610, \control_reg[7] , Stepper_Y_En_c, 
            Stepper_Y_Dir_c, Stepper_Y_M2_c_2, Stepper_Y_M1_c_1, \read_size[2] , 
            n14121, \steps_reg[24] , n32385, n32381, n32382, \steps_reg[20] , 
            n3666, n32383, \steps_reg[4] , \steps_reg[1] , \register_addr[1] , 
            fault_latched, VCC_net, GND_net, Stepper_Y_nFault_c, \read_size[0] , 
            n32, \register_addr[2] , \register_addr[3] , \register_addr[4] , 
            n28196, Stepper_Y_M0_c_0, n579, prev_step_clk, step_clk, 
            prev_select, n30374, read_value, n9128, n26485, \register_addr[0] , 
            n30370, n30380, n30421, \register_addr[5] , limit_c_1, 
            Stepper_Y_Step_c, n30489, n30491, \select[4] , n30427, 
            n30406, n30417, n28184, n32380, n30316, n13269, n30331, 
            rw, n22, n30311, n21533, n28324, n30479, n28323, n12, 
            n28172, n19585, n30342, \div_factor_reg[24] , n28672, 
            \div_factor_reg[1] , n49, \div_factor_reg[20] , n17, n8263) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n8894;
    input n32384;
    input [31:0]databus;
    input n608;
    input n610;
    output \control_reg[7] ;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output Stepper_Y_M2_c_2;
    output Stepper_Y_M1_c_1;
    output \read_size[2] ;
    input n14121;
    output \steps_reg[24] ;
    input n32385;
    input n32381;
    input n32382;
    output \steps_reg[20] ;
    input n3666;
    input n32383;
    output \steps_reg[4] ;
    output \steps_reg[1] ;
    input \register_addr[1] ;
    output fault_latched;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    output \read_size[0] ;
    input n32;
    input \register_addr[2] ;
    input \register_addr[3] ;
    input \register_addr[4] ;
    output n28196;
    output Stepper_Y_M0_c_0;
    input n579;
    output prev_step_clk;
    output step_clk;
    output prev_select;
    input n30374;
    output [31:0]read_value;
    input n9128;
    output n26485;
    input \register_addr[0] ;
    output n30370;
    output n30380;
    output n30421;
    input \register_addr[5] ;
    input limit_c_1;
    output Stepper_Y_Step_c;
    output n30489;
    input n30491;
    input \select[4] ;
    output n30427;
    output n30406;
    output n30417;
    output n28184;
    input n32380;
    input n30316;
    input n13269;
    input n30331;
    input rw;
    input n22;
    input n30311;
    input n21533;
    output n28324;
    input n30479;
    output n28323;
    input n12;
    output n28172;
    output n19585;
    input n30342;
    output \div_factor_reg[24] ;
    input n28672;
    output \div_factor_reg[1] ;
    input n49;
    output \div_factor_reg[20] ;
    input n17;
    input n8263;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n13318, n30309, n10718;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n13335, n28170;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n3667;
    wire [31:0]n224;
    
    wire n28637, n28322, n28638, limit_latched, n182, prev_limit_latched, 
        n28696, n49_c, n62, n58, n50, n41, n60, n54, n42, 
        n52, n38, n56, n46, n28639;
    wire [31:0]n100;
    
    wire n24, n30453, int_step, n25950, n25949, n25948, n25947, 
        n25946, n25945, n25944, n25943, n25942, n25941, n25940, 
        n25939, n29, n25938;
    wire [31:0]n99;
    
    wire n25937, n25936, n25935;
    wire [31:0]n6577;
    
    wire n28694, n28695, n19589;
    wire [7:0]n8262;
    wire [31:0]n6541;
    
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n8894), .PD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n8894), .PD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n8894), .PD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n8894), .PD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n8894), .PD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n8894), .PD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n8894), .PD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n13318), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n13318), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n30309), .CD(n10718), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n30309), .PD(n32384), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n30309), .PD(n32384), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n13335), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n30309), .PD(n32384), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n13335), .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n30309), .PD(n32384), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n28170), .SP(n14121), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3667[31]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3667[30]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3667[29]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3667[28]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3667[27]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3667[26]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3667[25]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3667[24]), .CK(debug_c_c), .CD(n32384), 
            .Q(\steps_reg[24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3667[23]), .CK(debug_c_c), .CD(n32385), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3667[22]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3667[21]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3667[20]), .CK(debug_c_c), .CD(n32382), 
            .Q(\steps_reg[20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3667[19]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3667[18]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3667[17]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    LUT4 mux_1514_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3666), 
         .Z(n3667[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i27_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i16 (.D(n3667[16]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3667[15]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3667[14]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3667[13]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3667[12]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3667[11]), .CK(debug_c_c), .CD(n32383), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3667[10]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3667[9]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3667[8]), .CK(debug_c_c), .CD(n32383), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3667[7]), .CK(debug_c_c), .CD(n32383), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3667[6]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3667[5]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3667[4]), .CK(debug_c_c), .CD(n32383), 
            .Q(\steps_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3667[3]), .CK(debug_c_c), .CD(n32383), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3667[2]), .CK(debug_c_c), .CD(n32383), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3667[1]), .CK(debug_c_c), .CD(n32383), 
            .Q(\steps_reg[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i21484_3_lut (.A(Stepper_Y_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n28637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21484_3_lut.init = 16'hcaca;
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3667[0]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n28322), .SP(n14121), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i21485_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n28638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21485_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .C(\register_addr[4] ), .Z(n28196)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    FD1P3AX control_reg_i1 (.D(n579), .SP(n13335), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13318), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n30374), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n28696), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i31_4_lut (.A(n49_c), .B(n62), .C(n58), .D(n50), .Z(n26485)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[16]), .Z(n49_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(steps_reg[9]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 equal_55_i8_1_lut_rep_361_2_lut_3_lut_4_lut (.A(\register_addr[2] ), 
         .B(\register_addr[3] ), .C(\register_addr[0] ), .D(\register_addr[1] ), 
         .Z(n30370)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_55_i8_1_lut_rep_361_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_371_3_lut_4_lut (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .C(\register_addr[0] ), .D(\register_addr[1] ), .Z(n30380)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_371_3_lut_4_lut.init = 16'hfffe;
    PFUMX i21486 (.BLUT(n28637), .ALUT(n28638), .C0(\register_addr[0] ), 
          .Z(n28639));
    LUT4 i22_4_lut (.A(steps_reg[2]), .B(\steps_reg[4] ), .C(\steps_reg[20] ), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(\steps_reg[1] ), 
         .D(steps_reg[3]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[6]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[8]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(\steps_reg[24] ), .B(steps_reg[0]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i14618_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14618_4_lut.init = 16'hc088;
    LUT4 i14619_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14619_4_lut.init = 16'hc088;
    LUT4 i14620_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14620_4_lut.init = 16'hc088;
    LUT4 i14621_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14621_4_lut.init = 16'hc088;
    LUT4 i14622_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14622_4_lut.init = 16'hc088;
    LUT4 i14623_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14623_4_lut.init = 16'hc088;
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[16]), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n24)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i14624_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14624_4_lut.init = 16'hc088;
    LUT4 i14625_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14625_4_lut.init = 16'hc088;
    LUT4 i14626_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14626_4_lut.init = 16'hc088;
    LUT4 i14627_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14627_4_lut.init = 16'hc088;
    LUT4 i14628_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14628_4_lut.init = 16'hc088;
    LUT4 i14629_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14629_4_lut.init = 16'hc088;
    LUT4 i14630_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14630_4_lut.init = 16'hc088;
    LUT4 mux_1514_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3666), .Z(n3667[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(n30421), .B(\register_addr[5] ), .C(\register_addr[4] ), 
         .Z(n28170)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i2_3_lut.init = 16'h2020;
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_444 (.A(\register_addr[5] ), .B(\register_addr[4] ), 
         .Z(n30453)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i1_2_lut_rep_444.init = 16'hbbbb;
    LUT4 mux_1514_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3666), 
         .Z(n3667[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3666), 
         .Z(n3667[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3666), 
         .Z(n3667[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3666), 
         .Z(n3667[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i29_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1514_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3666), 
         .Z(n3667[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i28_3_lut.init = 16'hcaca;
    LUT4 equal_1539_i11_2_lut_rep_480 (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .Z(n30489)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_1539_i11_2_lut_rep_480.init = 16'heeee;
    LUT4 i1_3_lut_rep_418_4_lut (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .C(n30491), .D(\select[4] ), .Z(n30427)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_3_lut_rep_418_4_lut.init = 16'h0100;
    LUT4 i14775_2_lut_rep_397_3_lut (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .C(\register_addr[1] ), .Z(n30406)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i14775_2_lut_rep_397_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_408_3_lut (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .C(\register_addr[5] ), .Z(n30417)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_408_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .C(\register_addr[4] ), .D(\register_addr[5] ), .Z(n28184)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i21701_2_lut_4_lut_4_lut (.A(n30453), .B(n32380), .C(n30316), 
         .D(n13269), .Z(n13335)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i21701_2_lut_4_lut_4_lut.init = 16'hccdc;
    LUT4 i21705_3_lut_rep_300_4_lut_4_lut (.A(n30453), .B(n13269), .C(n30331), 
         .D(rw), .Z(n30309)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i21705_3_lut_rep_300_4_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_201 (.A(n8894), .B(n32380), .Z(n13318)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_201.init = 16'heeee;
    LUT4 mux_1514_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3666), 
         .Z(n3667[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i26_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_412_4_lut (.A(\register_addr[2] ), .B(\register_addr[3] ), 
         .C(n30491), .D(\register_addr[1] ), .Z(n30421)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i2_3_lut_rep_412_4_lut.init = 16'h0100;
    FD1P3AX int_step_182 (.D(n30311), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i21661_2_lut_2_lut_3_lut_4_lut (.A(n30489), .B(\register_addr[1] ), 
         .C(n21533), .D(n30491), .Z(n28324)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21661_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i21664_2_lut_2_lut_3_lut_4_lut (.A(n30489), .B(\register_addr[1] ), 
         .C(n30479), .D(n30491), .Z(n28323)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21664_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i21667_2_lut_2_lut_3_lut_4_lut (.A(n30489), .B(\register_addr[1] ), 
         .C(n30453), .D(n30491), .Z(n28322)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21667_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n12), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n24), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n30489), .B(\register_addr[1] ), .C(n30491), 
         .D(n21533), .Z(n28172)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 mux_1514_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3666), 
         .Z(n3667[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i25_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    LUT4 mux_1514_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3666), 
         .Z(n3667[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3666), 
         .Z(n3667[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3666), 
         .Z(n3667[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3666), 
         .Z(n3667[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3666), 
         .Z(n3667[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3666), 
         .Z(n3667[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3666), 
         .Z(n3667[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3666), 
         .Z(n3667[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i17_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25950), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    LUT4 mux_1514_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3666), 
         .Z(n3667[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i16_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25949), .COUT(n25950), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25948), .COUT(n25949), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25947), .COUT(n25948), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25946), .COUT(n25947), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    LUT4 mux_1514_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3666), 
         .Z(n3667[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i15_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25945), .COUT(n25946), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25944), .COUT(n25945), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    LUT4 mux_1514_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3666), 
         .Z(n3667[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3666), 
         .Z(n3667[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i13_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25943), .COUT(n25944), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25942), .COUT(n25943), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25941), .COUT(n25942), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    LUT4 mux_1514_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3666), 
         .Z(n3667[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3666), 
         .Z(n3667[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3666), .Z(n3667[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3666), .Z(n3667[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3666), .Z(n3667[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3666), .Z(n3667[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i7_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25940), .COUT(n25941), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25939), .COUT(n25940), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_202 (.A(div_factor_reg[8]), .B(n19585), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_202.init = 16'hc088;
    LUT4 i1_2_lut_adj_203 (.A(\register_addr[1] ), .B(n9128), .Z(n19585)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_2_lut_adj_203.init = 16'h2222;
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25938), .COUT(n25939), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_204 (.A(n19585), .B(div_factor_reg[25]), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n99[25])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_204.init = 16'ha088;
    LUT4 i1_4_lut_adj_205 (.A(n19585), .B(div_factor_reg[26]), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n99[26])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_205.init = 16'ha088;
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25937), .COUT(n25938), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25936), .COUT(n25937), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_206 (.A(n19585), .B(div_factor_reg[27]), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n99[27])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_206.init = 16'ha088;
    LUT4 i1_4_lut_adj_207 (.A(n19585), .B(div_factor_reg[28]), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n99[28])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_207.init = 16'ha088;
    CCU2D sub_125_add_2_3 (.A0(\steps_reg[1] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25935), .COUT(n25936), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_208 (.A(n19585), .B(div_factor_reg[29]), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n99[29])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_208.init = 16'ha088;
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n25935), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_209 (.A(n19585), .B(div_factor_reg[30]), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n99[30])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_209.init = 16'ha088;
    LUT4 i14939_4_lut (.A(div_factor_reg[31]), .B(n19585), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n99[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i14939_4_lut.init = 16'hc088;
    LUT4 mux_1514_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3666), .Z(n3667[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3666), .Z(n3667[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3666), .Z(n3667[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i4_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(\div_factor_reg[24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    LUT4 mux_1514_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3666), .Z(n3667[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1514_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3666), .Z(n3667[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1514_i2_3_lut.init = 16'hcaca;
    LUT4 i4312_3_lut (.A(prev_limit_latched), .B(n32380), .C(limit_latched), 
         .Z(n10718)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i4312_3_lut.init = 16'hdcdc;
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n13318), .CD(n30342), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n28672), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n28639), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6577[3]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6577[4]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6577[5]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6577[6]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6577[7]), .SP(n14121), .CD(n9128), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(\div_factor_reg[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29), .SP(n14121), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n49), .SP(n14121), .CK(debug_c_c), .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n99[25]), .SP(n14121), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n99[26]), .SP(n14121), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n99[27]), .SP(n14121), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n99[28]), .SP(n14121), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n99[29]), .SP(n14121), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n99[30]), .SP(n14121), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n99[31]), .SP(n14121), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n13318), .CD(n32384), 
            .CK(debug_c_c), .Q(\div_factor_reg[20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    LUT4 i21541_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n28694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21541_3_lut.init = 16'hcaca;
    LUT4 i21542_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n28695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21542_3_lut.init = 16'hcaca;
    LUT4 i13198_3_lut (.A(control_reg[4]), .B(div_factor_reg[4]), .C(\register_addr[1] ), 
         .Z(n19589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13198_3_lut.init = 16'hcaca;
    LUT4 i14636_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8262[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14636_2_lut.init = 16'h2222;
    LUT4 mux_1915_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n6541[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1915_i4_3_lut.init = 16'hcaca;
    LUT4 i14635_2_lut (.A(Stepper_Y_Dir_c), .B(\register_addr[0] ), .Z(n8262[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14635_2_lut.init = 16'h2222;
    LUT4 mux_1915_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n6541[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1915_i6_3_lut.init = 16'hcaca;
    LUT4 i14634_2_lut (.A(Stepper_Y_En_c), .B(\register_addr[0] ), .Z(n8262[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14634_2_lut.init = 16'h2222;
    LUT4 mux_1915_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n6541[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1915_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1915_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6541[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1915_i8_3_lut.init = 16'hcaca;
    PFUMX i21543 (.BLUT(n28694), .ALUT(n28695), .C0(\register_addr[1] ), 
          .Z(n28696));
    PFUMX i13200 (.BLUT(n19589), .ALUT(n17), .C0(\register_addr[0] ), 
          .Z(n6577[4]));
    PFUMX mux_1919_i4 (.BLUT(n8262[3]), .ALUT(n6541[3]), .C0(\register_addr[1] ), 
          .Z(n6577[3]));
    PFUMX mux_1919_i6 (.BLUT(n8262[5]), .ALUT(n6541[5]), .C0(\register_addr[1] ), 
          .Z(n6577[5]));
    PFUMX mux_1919_i7 (.BLUT(n8262[6]), .ALUT(n6541[6]), .C0(\register_addr[1] ), 
          .Z(n6577[6]));
    PFUMX mux_1919_i8 (.BLUT(n8263), .ALUT(n6541[7]), .C0(\register_addr[1] ), 
          .Z(n6577[7]));
    ClockDivider_U7 step_clk_gen (.GND_net(GND_net), .n32380(n32380), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n32385(n32385), .div_factor_reg({div_factor_reg[31:25], 
            \div_factor_reg[24] , div_factor_reg[23:21], \div_factor_reg[20] , 
            div_factor_reg[19:2], \div_factor_reg[1] , div_factor_reg[0]})) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (GND_net, n32380, step_clk, debug_c_c, n32385, 
            div_factor_reg) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n32380;
    output step_clk;
    input debug_c_c;
    input n32385;
    input [31:0]div_factor_reg;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25884;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n25885, n25883, n25882, n25881, n25880, n25879, n25878, 
        n25877, n7782, n30302, n7816, n16213, n25876, n25875, 
        n25874, n25873, n25750;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n7747, n25872, n25749, n25748, n25871, n25747, n25746, 
        n25745, n25744, n25743, n25742, n25741, n25740, n25739, 
        n25738;
    wire [31:0]n134;
    
    wire n25737, n25736, n25735, n25734, n25733, n25732, n25731, 
        n25730, n25729, n25728, n25727, n25726, n25725, n25724, 
        n25723, n25722, n25721, n25720, n25719, n25990, n25718, 
        n25989, n25717, n25716, n25988, n25987, n25715, n25714, 
        n25986, n25713, n25712, n25985, n25711, n25710, n25984, 
        n25709, n25708, n25983, n25707, n25706, n25982, n25705, 
        n25704, n25981, n25703, n25980, n25979, n25978, n25977, 
        n25976, n25975, n25886;
    
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25884), .COUT(n25885), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25883), .COUT(n25884), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25882), .COUT(n25883), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25881), .COUT(n25882), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25880), .COUT(n25881), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25879), .COUT(n25880), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25878), .COUT(n25879), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25877), .COUT(n25878), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    LUT4 i1013_2_lut_rep_293 (.A(n7782), .B(n32380), .Z(n30302)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1013_2_lut_rep_293.init = 16'heeee;
    LUT4 i9801_2_lut_3_lut (.A(n7782), .B(n32380), .C(n7816), .Z(n16213)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9801_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25876), .COUT(n25877), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25875), .COUT(n25876), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25874), .COUT(n25875), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25873), .COUT(n25874), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25750), .S1(n7747));
    defparam sub_2019_add_2_33.INIT0 = 16'h5555;
    defparam sub_2019_add_2_33.INIT1 = 16'h0000;
    defparam sub_2019_add_2_33.INJECT1_0 = "NO";
    defparam sub_2019_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25872), .COUT(n25873), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25749), .COUT(n25750));
    defparam sub_2019_add_2_31.INIT0 = 16'h5999;
    defparam sub_2019_add_2_31.INIT1 = 16'h5999;
    defparam sub_2019_add_2_31.INJECT1_0 = "NO";
    defparam sub_2019_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25748), .COUT(n25749));
    defparam sub_2019_add_2_29.INIT0 = 16'h5999;
    defparam sub_2019_add_2_29.INIT1 = 16'h5999;
    defparam sub_2019_add_2_29.INJECT1_0 = "NO";
    defparam sub_2019_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25871), .COUT(n25872), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25871), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25747), .COUT(n25748));
    defparam sub_2019_add_2_27.INIT0 = 16'h5999;
    defparam sub_2019_add_2_27.INIT1 = 16'h5999;
    defparam sub_2019_add_2_27.INJECT1_0 = "NO";
    defparam sub_2019_add_2_27.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7747), .CK(debug_c_c), .CD(n32385), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2019_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25746), .COUT(n25747));
    defparam sub_2019_add_2_25.INIT0 = 16'h5999;
    defparam sub_2019_add_2_25.INIT1 = 16'h5999;
    defparam sub_2019_add_2_25.INJECT1_0 = "NO";
    defparam sub_2019_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25745), .COUT(n25746));
    defparam sub_2019_add_2_23.INIT0 = 16'h5999;
    defparam sub_2019_add_2_23.INIT1 = 16'h5999;
    defparam sub_2019_add_2_23.INJECT1_0 = "NO";
    defparam sub_2019_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25744), .COUT(n25745));
    defparam sub_2019_add_2_21.INIT0 = 16'h5999;
    defparam sub_2019_add_2_21.INIT1 = 16'h5999;
    defparam sub_2019_add_2_21.INJECT1_0 = "NO";
    defparam sub_2019_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25743), .COUT(n25744));
    defparam sub_2019_add_2_19.INIT0 = 16'h5999;
    defparam sub_2019_add_2_19.INIT1 = 16'h5999;
    defparam sub_2019_add_2_19.INJECT1_0 = "NO";
    defparam sub_2019_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25742), .COUT(n25743));
    defparam sub_2019_add_2_17.INIT0 = 16'h5999;
    defparam sub_2019_add_2_17.INIT1 = 16'h5999;
    defparam sub_2019_add_2_17.INJECT1_0 = "NO";
    defparam sub_2019_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25741), .COUT(n25742));
    defparam sub_2019_add_2_15.INIT0 = 16'h5999;
    defparam sub_2019_add_2_15.INIT1 = 16'h5999;
    defparam sub_2019_add_2_15.INJECT1_0 = "NO";
    defparam sub_2019_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25740), .COUT(n25741));
    defparam sub_2019_add_2_13.INIT0 = 16'h5999;
    defparam sub_2019_add_2_13.INIT1 = 16'h5999;
    defparam sub_2019_add_2_13.INJECT1_0 = "NO";
    defparam sub_2019_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25739), .COUT(n25740));
    defparam sub_2019_add_2_11.INIT0 = 16'h5999;
    defparam sub_2019_add_2_11.INIT1 = 16'h5999;
    defparam sub_2019_add_2_11.INJECT1_0 = "NO";
    defparam sub_2019_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25738), .COUT(n25739));
    defparam sub_2019_add_2_9.INIT0 = 16'h5999;
    defparam sub_2019_add_2_9.INIT1 = 16'h5999;
    defparam sub_2019_add_2_9.INJECT1_0 = "NO";
    defparam sub_2019_add_2_9.INJECT1_1 = "NO";
    FD1S3IX count_2612__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i0.GSR = "ENABLED";
    CCU2D sub_2019_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25737), .COUT(n25738));
    defparam sub_2019_add_2_7.INIT0 = 16'h5999;
    defparam sub_2019_add_2_7.INIT1 = 16'h5999;
    defparam sub_2019_add_2_7.INJECT1_0 = "NO";
    defparam sub_2019_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25736), .COUT(n25737));
    defparam sub_2019_add_2_5.INIT0 = 16'h5999;
    defparam sub_2019_add_2_5.INIT1 = 16'h5999;
    defparam sub_2019_add_2_5.INJECT1_0 = "NO";
    defparam sub_2019_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25735), .COUT(n25736));
    defparam sub_2019_add_2_3.INIT0 = 16'h5999;
    defparam sub_2019_add_2_3.INIT1 = 16'h5999;
    defparam sub_2019_add_2_3.INJECT1_0 = "NO";
    defparam sub_2019_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2019_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n25735));
    defparam sub_2019_add_2_1.INIT0 = 16'h0000;
    defparam sub_2019_add_2_1.INIT1 = 16'h5999;
    defparam sub_2019_add_2_1.INJECT1_0 = "NO";
    defparam sub_2019_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25734), .S1(n7782));
    defparam sub_2021_add_2_33.INIT0 = 16'h5999;
    defparam sub_2021_add_2_33.INIT1 = 16'h0000;
    defparam sub_2021_add_2_33.INJECT1_0 = "NO";
    defparam sub_2021_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25733), .COUT(n25734));
    defparam sub_2021_add_2_31.INIT0 = 16'h5999;
    defparam sub_2021_add_2_31.INIT1 = 16'h5999;
    defparam sub_2021_add_2_31.INJECT1_0 = "NO";
    defparam sub_2021_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25732), .COUT(n25733));
    defparam sub_2021_add_2_29.INIT0 = 16'h5999;
    defparam sub_2021_add_2_29.INIT1 = 16'h5999;
    defparam sub_2021_add_2_29.INJECT1_0 = "NO";
    defparam sub_2021_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25731), .COUT(n25732));
    defparam sub_2021_add_2_27.INIT0 = 16'h5999;
    defparam sub_2021_add_2_27.INIT1 = 16'h5999;
    defparam sub_2021_add_2_27.INJECT1_0 = "NO";
    defparam sub_2021_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25730), .COUT(n25731));
    defparam sub_2021_add_2_25.INIT0 = 16'h5999;
    defparam sub_2021_add_2_25.INIT1 = 16'h5999;
    defparam sub_2021_add_2_25.INJECT1_0 = "NO";
    defparam sub_2021_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25729), .COUT(n25730));
    defparam sub_2021_add_2_23.INIT0 = 16'h5999;
    defparam sub_2021_add_2_23.INIT1 = 16'h5999;
    defparam sub_2021_add_2_23.INJECT1_0 = "NO";
    defparam sub_2021_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25728), .COUT(n25729));
    defparam sub_2021_add_2_21.INIT0 = 16'h5999;
    defparam sub_2021_add_2_21.INIT1 = 16'h5999;
    defparam sub_2021_add_2_21.INJECT1_0 = "NO";
    defparam sub_2021_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25727), .COUT(n25728));
    defparam sub_2021_add_2_19.INIT0 = 16'h5999;
    defparam sub_2021_add_2_19.INIT1 = 16'h5999;
    defparam sub_2021_add_2_19.INJECT1_0 = "NO";
    defparam sub_2021_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25726), .COUT(n25727));
    defparam sub_2021_add_2_17.INIT0 = 16'h5999;
    defparam sub_2021_add_2_17.INIT1 = 16'h5999;
    defparam sub_2021_add_2_17.INJECT1_0 = "NO";
    defparam sub_2021_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25725), .COUT(n25726));
    defparam sub_2021_add_2_15.INIT0 = 16'h5999;
    defparam sub_2021_add_2_15.INIT1 = 16'h5999;
    defparam sub_2021_add_2_15.INJECT1_0 = "NO";
    defparam sub_2021_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25724), .COUT(n25725));
    defparam sub_2021_add_2_13.INIT0 = 16'h5999;
    defparam sub_2021_add_2_13.INIT1 = 16'h5999;
    defparam sub_2021_add_2_13.INJECT1_0 = "NO";
    defparam sub_2021_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25723), .COUT(n25724));
    defparam sub_2021_add_2_11.INIT0 = 16'h5999;
    defparam sub_2021_add_2_11.INIT1 = 16'h5999;
    defparam sub_2021_add_2_11.INJECT1_0 = "NO";
    defparam sub_2021_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25722), .COUT(n25723));
    defparam sub_2021_add_2_9.INIT0 = 16'h5999;
    defparam sub_2021_add_2_9.INIT1 = 16'h5999;
    defparam sub_2021_add_2_9.INJECT1_0 = "NO";
    defparam sub_2021_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25721), .COUT(n25722));
    defparam sub_2021_add_2_7.INIT0 = 16'h5999;
    defparam sub_2021_add_2_7.INIT1 = 16'h5999;
    defparam sub_2021_add_2_7.INJECT1_0 = "NO";
    defparam sub_2021_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25720), .COUT(n25721));
    defparam sub_2021_add_2_5.INIT0 = 16'h5999;
    defparam sub_2021_add_2_5.INIT1 = 16'h5999;
    defparam sub_2021_add_2_5.INJECT1_0 = "NO";
    defparam sub_2021_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25719), .COUT(n25720));
    defparam sub_2021_add_2_3.INIT0 = 16'h5999;
    defparam sub_2021_add_2_3.INIT1 = 16'h5999;
    defparam sub_2021_add_2_3.INJECT1_0 = "NO";
    defparam sub_2021_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25990), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_33.INIT1 = 16'h0000;
    defparam count_2612_add_4_33.INJECT1_0 = "NO";
    defparam count_2612_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_2021_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n25719));
    defparam sub_2021_add_2_1.INIT0 = 16'h0000;
    defparam sub_2021_add_2_1.INIT1 = 16'h5999;
    defparam sub_2021_add_2_1.INJECT1_0 = "NO";
    defparam sub_2021_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25718), .S1(n7816));
    defparam sub_2022_add_2_33.INIT0 = 16'hf555;
    defparam sub_2022_add_2_33.INIT1 = 16'h0000;
    defparam sub_2022_add_2_33.INJECT1_0 = "NO";
    defparam sub_2022_add_2_33.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25989), .COUT(n25990), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_31.INJECT1_0 = "NO";
    defparam count_2612_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25717), .COUT(n25718));
    defparam sub_2022_add_2_31.INIT0 = 16'hf555;
    defparam sub_2022_add_2_31.INIT1 = 16'hf555;
    defparam sub_2022_add_2_31.INJECT1_0 = "NO";
    defparam sub_2022_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25716), .COUT(n25717));
    defparam sub_2022_add_2_29.INIT0 = 16'hf555;
    defparam sub_2022_add_2_29.INIT1 = 16'hf555;
    defparam sub_2022_add_2_29.INJECT1_0 = "NO";
    defparam sub_2022_add_2_29.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25988), .COUT(n25989), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_29.INJECT1_0 = "NO";
    defparam count_2612_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25987), .COUT(n25988), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_27.INJECT1_0 = "NO";
    defparam count_2612_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25715), .COUT(n25716));
    defparam sub_2022_add_2_27.INIT0 = 16'hf555;
    defparam sub_2022_add_2_27.INIT1 = 16'hf555;
    defparam sub_2022_add_2_27.INJECT1_0 = "NO";
    defparam sub_2022_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25714), .COUT(n25715));
    defparam sub_2022_add_2_25.INIT0 = 16'hf555;
    defparam sub_2022_add_2_25.INIT1 = 16'hf555;
    defparam sub_2022_add_2_25.INJECT1_0 = "NO";
    defparam sub_2022_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25986), .COUT(n25987), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_25.INJECT1_0 = "NO";
    defparam count_2612_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25713), .COUT(n25714));
    defparam sub_2022_add_2_23.INIT0 = 16'hf555;
    defparam sub_2022_add_2_23.INIT1 = 16'hf555;
    defparam sub_2022_add_2_23.INJECT1_0 = "NO";
    defparam sub_2022_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25712), .COUT(n25713));
    defparam sub_2022_add_2_21.INIT0 = 16'hf555;
    defparam sub_2022_add_2_21.INIT1 = 16'hf555;
    defparam sub_2022_add_2_21.INJECT1_0 = "NO";
    defparam sub_2022_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25985), .COUT(n25986), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_23.INJECT1_0 = "NO";
    defparam count_2612_add_4_23.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25711), .COUT(n25712));
    defparam sub_2022_add_2_19.INIT0 = 16'hf555;
    defparam sub_2022_add_2_19.INIT1 = 16'hf555;
    defparam sub_2022_add_2_19.INJECT1_0 = "NO";
    defparam sub_2022_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25710), .COUT(n25711));
    defparam sub_2022_add_2_17.INIT0 = 16'hf555;
    defparam sub_2022_add_2_17.INIT1 = 16'hf555;
    defparam sub_2022_add_2_17.INJECT1_0 = "NO";
    defparam sub_2022_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25984), .COUT(n25985), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_21.INJECT1_0 = "NO";
    defparam count_2612_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25709), .COUT(n25710));
    defparam sub_2022_add_2_15.INIT0 = 16'hf555;
    defparam sub_2022_add_2_15.INIT1 = 16'hf555;
    defparam sub_2022_add_2_15.INJECT1_0 = "NO";
    defparam sub_2022_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25708), .COUT(n25709));
    defparam sub_2022_add_2_13.INIT0 = 16'hf555;
    defparam sub_2022_add_2_13.INIT1 = 16'hf555;
    defparam sub_2022_add_2_13.INJECT1_0 = "NO";
    defparam sub_2022_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25983), .COUT(n25984), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_19.INJECT1_0 = "NO";
    defparam count_2612_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25707), .COUT(n25708));
    defparam sub_2022_add_2_11.INIT0 = 16'hf555;
    defparam sub_2022_add_2_11.INIT1 = 16'hf555;
    defparam sub_2022_add_2_11.INJECT1_0 = "NO";
    defparam sub_2022_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25706), .COUT(n25707));
    defparam sub_2022_add_2_9.INIT0 = 16'hf555;
    defparam sub_2022_add_2_9.INIT1 = 16'hf555;
    defparam sub_2022_add_2_9.INJECT1_0 = "NO";
    defparam sub_2022_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25982), .COUT(n25983), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_17.INJECT1_0 = "NO";
    defparam count_2612_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25705), .COUT(n25706));
    defparam sub_2022_add_2_7.INIT0 = 16'hf555;
    defparam sub_2022_add_2_7.INIT1 = 16'hf555;
    defparam sub_2022_add_2_7.INJECT1_0 = "NO";
    defparam sub_2022_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25704), .COUT(n25705));
    defparam sub_2022_add_2_5.INIT0 = 16'hf555;
    defparam sub_2022_add_2_5.INIT1 = 16'hf555;
    defparam sub_2022_add_2_5.INJECT1_0 = "NO";
    defparam sub_2022_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25981), .COUT(n25982), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_15.INJECT1_0 = "NO";
    defparam count_2612_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25703), .COUT(n25704));
    defparam sub_2022_add_2_3.INIT0 = 16'hf555;
    defparam sub_2022_add_2_3.INIT1 = 16'hf555;
    defparam sub_2022_add_2_3.INJECT1_0 = "NO";
    defparam sub_2022_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25980), .COUT(n25981), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_13.INJECT1_0 = "NO";
    defparam count_2612_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25979), .COUT(n25980), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_11.INJECT1_0 = "NO";
    defparam count_2612_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_2022_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n25703));
    defparam sub_2022_add_2_1.INIT0 = 16'h0000;
    defparam sub_2022_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2022_add_2_1.INJECT1_0 = "NO";
    defparam sub_2022_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25978), .COUT(n25979), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_9.INJECT1_0 = "NO";
    defparam count_2612_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25977), .COUT(n25978), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_7.INJECT1_0 = "NO";
    defparam count_2612_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25976), .COUT(n25977), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_5.INJECT1_0 = "NO";
    defparam count_2612_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25975), .COUT(n25976), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2612_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2612_add_4_3.INJECT1_0 = "NO";
    defparam count_2612_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2612_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25975), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612_add_4_1.INIT0 = 16'hF000;
    defparam count_2612_add_4_1.INIT1 = 16'h0555;
    defparam count_2612_add_4_1.INJECT1_0 = "NO";
    defparam count_2612_add_4_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n30302), .PD(n16213), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1S3IX count_2612__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i1.GSR = "ENABLED";
    FD1S3IX count_2612__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i2.GSR = "ENABLED";
    FD1S3IX count_2612__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i3.GSR = "ENABLED";
    FD1S3IX count_2612__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i4.GSR = "ENABLED";
    FD1S3IX count_2612__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i5.GSR = "ENABLED";
    FD1S3IX count_2612__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i6.GSR = "ENABLED";
    FD1S3IX count_2612__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i7.GSR = "ENABLED";
    FD1S3IX count_2612__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i8.GSR = "ENABLED";
    FD1S3IX count_2612__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i9.GSR = "ENABLED";
    FD1S3IX count_2612__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i10.GSR = "ENABLED";
    FD1S3IX count_2612__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i11.GSR = "ENABLED";
    FD1S3IX count_2612__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i12.GSR = "ENABLED";
    FD1S3IX count_2612__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i13.GSR = "ENABLED";
    FD1S3IX count_2612__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i14.GSR = "ENABLED";
    FD1S3IX count_2612__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i15.GSR = "ENABLED";
    FD1S3IX count_2612__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i16.GSR = "ENABLED";
    FD1S3IX count_2612__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i17.GSR = "ENABLED";
    FD1S3IX count_2612__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i18.GSR = "ENABLED";
    FD1S3IX count_2612__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i19.GSR = "ENABLED";
    FD1S3IX count_2612__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i20.GSR = "ENABLED";
    FD1S3IX count_2612__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i21.GSR = "ENABLED";
    FD1S3IX count_2612__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i22.GSR = "ENABLED";
    FD1S3IX count_2612__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i23.GSR = "ENABLED";
    FD1S3IX count_2612__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i24.GSR = "ENABLED";
    FD1S3IX count_2612__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i25.GSR = "ENABLED";
    FD1S3IX count_2612__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i26.GSR = "ENABLED";
    FD1S3IX count_2612__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i27.GSR = "ENABLED";
    FD1S3IX count_2612__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i28.GSR = "ENABLED";
    FD1S3IX count_2612__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i29.GSR = "ENABLED";
    FD1S3IX count_2612__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i30.GSR = "ENABLED";
    FD1S3IX count_2612__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n30302), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2612__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n30302), .CD(n16213), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25886), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25885), .COUT(n25886), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (debug_c_c, n241, n32380, n7504, n30303, n28775, 
            n26601, n28723, n26592, GND_net, n28725, n26596, n28910, 
            n13624, n28859, n14284, n28857, n14306, n28855, n14307, 
            n28853, n14308, n28851, n14309, n28765, n26618, n28770, 
            n26607, n28773, n26604) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n241;
    input n32380;
    output n7504;
    output n30303;
    input n28775;
    output n26601;
    input n28723;
    output n26592;
    input GND_net;
    input n28725;
    output n26596;
    input n28910;
    output n13624;
    input n28859;
    output n14284;
    input n28857;
    output n14306;
    input n28855;
    output n14307;
    input n28853;
    output n14308;
    input n28851;
    output n14309;
    input n28765;
    output n26618;
    input n28770;
    output n26607;
    input n28773;
    output n26604;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire clk_255kHz, n26182, n7539, n26181;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n26180, n26179, n26178, n26177, n26176, n26175, n26174, 
        n26173, n26172, n26171, n26170, n2639;
    wire [31:0]n134;
    
    wire n26169, n26168, n26167, n26006, n26005, n26004, n26003, 
        n26002, n26001, n26000, n25999, n25998, n25997, n25996, 
        n25995, n25994, n25993, n25992, n25991, n26246, n26245, 
        n26244, n26243, n26242, n26241, n26240, n26239, n26238, 
        n26237, n26236, n26235, n26234, n26233, n26232;
    
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=518, LSE_RLINE=521 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_294 (.A(n32380), .B(clk_255kHz), .C(n7504), .Z(n30303)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_3_lut_rep_294.init = 16'h1010;
    LUT4 i21724_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28775), 
         .Z(n26601)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21724_2_lut_4_lut.init = 16'h1000;
    LUT4 i21672_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28723), 
         .Z(n26592)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21672_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_2009_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26182), .S0(n7539));
    defparam sub_2009_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2009_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2009_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2009_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26181), .COUT(n26182));
    defparam sub_2009_add_2_32.INIT0 = 16'h5555;
    defparam sub_2009_add_2_32.INIT1 = 16'h5555;
    defparam sub_2009_add_2_32.INJECT1_0 = "NO";
    defparam sub_2009_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26180), .COUT(n26181));
    defparam sub_2009_add_2_30.INIT0 = 16'h5555;
    defparam sub_2009_add_2_30.INIT1 = 16'h5555;
    defparam sub_2009_add_2_30.INJECT1_0 = "NO";
    defparam sub_2009_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26179), .COUT(n26180));
    defparam sub_2009_add_2_28.INIT0 = 16'h5555;
    defparam sub_2009_add_2_28.INIT1 = 16'h5555;
    defparam sub_2009_add_2_28.INJECT1_0 = "NO";
    defparam sub_2009_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26178), .COUT(n26179));
    defparam sub_2009_add_2_26.INIT0 = 16'h5555;
    defparam sub_2009_add_2_26.INIT1 = 16'h5555;
    defparam sub_2009_add_2_26.INJECT1_0 = "NO";
    defparam sub_2009_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26177), .COUT(n26178));
    defparam sub_2009_add_2_24.INIT0 = 16'h5555;
    defparam sub_2009_add_2_24.INIT1 = 16'h5555;
    defparam sub_2009_add_2_24.INJECT1_0 = "NO";
    defparam sub_2009_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26176), .COUT(n26177));
    defparam sub_2009_add_2_22.INIT0 = 16'h5555;
    defparam sub_2009_add_2_22.INIT1 = 16'h5555;
    defparam sub_2009_add_2_22.INJECT1_0 = "NO";
    defparam sub_2009_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26175), .COUT(n26176));
    defparam sub_2009_add_2_20.INIT0 = 16'h5555;
    defparam sub_2009_add_2_20.INIT1 = 16'h5555;
    defparam sub_2009_add_2_20.INJECT1_0 = "NO";
    defparam sub_2009_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26174), .COUT(n26175));
    defparam sub_2009_add_2_18.INIT0 = 16'h5555;
    defparam sub_2009_add_2_18.INIT1 = 16'h5555;
    defparam sub_2009_add_2_18.INJECT1_0 = "NO";
    defparam sub_2009_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26173), .COUT(n26174));
    defparam sub_2009_add_2_16.INIT0 = 16'h5555;
    defparam sub_2009_add_2_16.INIT1 = 16'h5555;
    defparam sub_2009_add_2_16.INJECT1_0 = "NO";
    defparam sub_2009_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26172), .COUT(n26173));
    defparam sub_2009_add_2_14.INIT0 = 16'h5555;
    defparam sub_2009_add_2_14.INIT1 = 16'h5555;
    defparam sub_2009_add_2_14.INJECT1_0 = "NO";
    defparam sub_2009_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26171), .COUT(n26172));
    defparam sub_2009_add_2_12.INIT0 = 16'h5555;
    defparam sub_2009_add_2_12.INIT1 = 16'h5555;
    defparam sub_2009_add_2_12.INJECT1_0 = "NO";
    defparam sub_2009_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26170), .COUT(n26171));
    defparam sub_2009_add_2_10.INIT0 = 16'h5555;
    defparam sub_2009_add_2_10.INIT1 = 16'h5555;
    defparam sub_2009_add_2_10.INJECT1_0 = "NO";
    defparam sub_2009_add_2_10.INJECT1_1 = "NO";
    FD1S3IX count_2608__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2639), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i0.GSR = "ENABLED";
    CCU2D sub_2009_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26169), .COUT(n26170));
    defparam sub_2009_add_2_8.INIT0 = 16'h5555;
    defparam sub_2009_add_2_8.INIT1 = 16'h5555;
    defparam sub_2009_add_2_8.INJECT1_0 = "NO";
    defparam sub_2009_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26168), .COUT(n26169));
    defparam sub_2009_add_2_6.INIT0 = 16'h5555;
    defparam sub_2009_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_2009_add_2_6.INJECT1_0 = "NO";
    defparam sub_2009_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26167), .COUT(n26168));
    defparam sub_2009_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2009_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_2009_add_2_4.INJECT1_0 = "NO";
    defparam sub_2009_add_2_4.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26006), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_33.INIT1 = 16'h0000;
    defparam count_2608_add_4_33.INJECT1_0 = "NO";
    defparam count_2608_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26005), .COUT(n26006), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_31.INJECT1_0 = "NO";
    defparam count_2608_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26004), .COUT(n26005), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_29.INJECT1_0 = "NO";
    defparam count_2608_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26167));
    defparam sub_2009_add_2_2.INIT0 = 16'h0000;
    defparam sub_2009_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2009_add_2_2.INJECT1_0 = "NO";
    defparam sub_2009_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26003), .COUT(n26004), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_27.INJECT1_0 = "NO";
    defparam count_2608_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26002), .COUT(n26003), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_25.INJECT1_0 = "NO";
    defparam count_2608_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26001), .COUT(n26002), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_23.INJECT1_0 = "NO";
    defparam count_2608_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26000), .COUT(n26001), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_21.INJECT1_0 = "NO";
    defparam count_2608_add_4_21.INJECT1_1 = "NO";
    LUT4 i21674_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28725), 
         .Z(n26596)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21674_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2608_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25999), .COUT(n26000), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_19.INJECT1_0 = "NO";
    defparam count_2608_add_4_19.INJECT1_1 = "NO";
    LUT4 i21859_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28910), 
         .Z(n13624)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21859_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2608_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25998), .COUT(n25999), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_17.INJECT1_0 = "NO";
    defparam count_2608_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25997), .COUT(n25998), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_15.INJECT1_0 = "NO";
    defparam count_2608_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25996), .COUT(n25997), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_13.INJECT1_0 = "NO";
    defparam count_2608_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25995), .COUT(n25996), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_11.INJECT1_0 = "NO";
    defparam count_2608_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25994), .COUT(n25995), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_9.INJECT1_0 = "NO";
    defparam count_2608_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25993), .COUT(n25994), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_7.INJECT1_0 = "NO";
    defparam count_2608_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25992), .COUT(n25993), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_5.INJECT1_0 = "NO";
    defparam count_2608_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25991), .COUT(n25992), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2608_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2608_add_4_3.INJECT1_0 = "NO";
    defparam count_2608_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2608_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25991), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608_add_4_1.INIT0 = 16'hF000;
    defparam count_2608_add_4_1.INIT1 = 16'h0555;
    defparam count_2608_add_4_1.INJECT1_0 = "NO";
    defparam count_2608_add_4_1.INJECT1_1 = "NO";
    LUT4 i21808_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28859), 
         .Z(n14284)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21808_2_lut_4_lut.init = 16'h1000;
    LUT4 i21806_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28857), 
         .Z(n14306)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21806_2_lut_4_lut.init = 16'h1000;
    LUT4 i956_2_lut (.A(n7539), .B(n32380), .Z(n2639)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i956_2_lut.init = 16'heeee;
    LUT4 i21804_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28855), 
         .Z(n14307)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21804_2_lut_4_lut.init = 16'h1000;
    LUT4 i21802_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28853), 
         .Z(n14308)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21802_2_lut_4_lut.init = 16'h1000;
    LUT4 i21800_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28851), 
         .Z(n14309)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21800_2_lut_4_lut.init = 16'h1000;
    FD1S3IX count_2608__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2639), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i1.GSR = "ENABLED";
    FD1S3IX count_2608__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2639), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i2.GSR = "ENABLED";
    FD1S3IX count_2608__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2639), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i3.GSR = "ENABLED";
    FD1S3IX count_2608__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2639), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i4.GSR = "ENABLED";
    FD1S3IX count_2608__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2639), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i5.GSR = "ENABLED";
    FD1S3IX count_2608__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2639), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i6.GSR = "ENABLED";
    FD1S3IX count_2608__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2639), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i7.GSR = "ENABLED";
    FD1S3IX count_2608__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2639), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i8.GSR = "ENABLED";
    FD1S3IX count_2608__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2639), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i9.GSR = "ENABLED";
    FD1S3IX count_2608__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i10.GSR = "ENABLED";
    FD1S3IX count_2608__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i11.GSR = "ENABLED";
    FD1S3IX count_2608__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i12.GSR = "ENABLED";
    FD1S3IX count_2608__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i13.GSR = "ENABLED";
    FD1S3IX count_2608__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i14.GSR = "ENABLED";
    FD1S3IX count_2608__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i15.GSR = "ENABLED";
    FD1S3IX count_2608__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i16.GSR = "ENABLED";
    FD1S3IX count_2608__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i17.GSR = "ENABLED";
    FD1S3IX count_2608__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i18.GSR = "ENABLED";
    FD1S3IX count_2608__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i19.GSR = "ENABLED";
    FD1S3IX count_2608__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i20.GSR = "ENABLED";
    FD1S3IX count_2608__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i21.GSR = "ENABLED";
    FD1S3IX count_2608__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i22.GSR = "ENABLED";
    FD1S3IX count_2608__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i23.GSR = "ENABLED";
    FD1S3IX count_2608__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i24.GSR = "ENABLED";
    FD1S3IX count_2608__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i25.GSR = "ENABLED";
    FD1S3IX count_2608__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i26.GSR = "ENABLED";
    FD1S3IX count_2608__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i27.GSR = "ENABLED";
    FD1S3IX count_2608__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i28.GSR = "ENABLED";
    FD1S3IX count_2608__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i29.GSR = "ENABLED";
    FD1S3IX count_2608__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i30.GSR = "ENABLED";
    FD1S3IX count_2608__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2639), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2608__i31.GSR = "ENABLED";
    LUT4 i21714_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28765), 
         .Z(n26618)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21714_2_lut_4_lut.init = 16'h1000;
    LUT4 i21719_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28770), 
         .Z(n26607)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21719_2_lut_4_lut.init = 16'h1000;
    LUT4 i21722_2_lut_4_lut (.A(n32380), .B(clk_255kHz), .C(n7504), .D(n28773), 
         .Z(n26604)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21722_2_lut_4_lut.init = 16'h1000;
    CCU2D add_19120_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26246), 
          .S1(n7504));
    defparam add_19120_32.INIT0 = 16'h5555;
    defparam add_19120_32.INIT1 = 16'h0000;
    defparam add_19120_32.INJECT1_0 = "NO";
    defparam add_19120_32.INJECT1_1 = "NO";
    CCU2D add_19120_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26245), .COUT(n26246));
    defparam add_19120_30.INIT0 = 16'h5555;
    defparam add_19120_30.INIT1 = 16'h5555;
    defparam add_19120_30.INJECT1_0 = "NO";
    defparam add_19120_30.INJECT1_1 = "NO";
    CCU2D add_19120_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26244), .COUT(n26245));
    defparam add_19120_28.INIT0 = 16'h5555;
    defparam add_19120_28.INIT1 = 16'h5555;
    defparam add_19120_28.INJECT1_0 = "NO";
    defparam add_19120_28.INJECT1_1 = "NO";
    CCU2D add_19120_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26243), .COUT(n26244));
    defparam add_19120_26.INIT0 = 16'h5555;
    defparam add_19120_26.INIT1 = 16'h5555;
    defparam add_19120_26.INJECT1_0 = "NO";
    defparam add_19120_26.INJECT1_1 = "NO";
    CCU2D add_19120_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26242), .COUT(n26243));
    defparam add_19120_24.INIT0 = 16'h5555;
    defparam add_19120_24.INIT1 = 16'h5555;
    defparam add_19120_24.INJECT1_0 = "NO";
    defparam add_19120_24.INJECT1_1 = "NO";
    CCU2D add_19120_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26241), .COUT(n26242));
    defparam add_19120_22.INIT0 = 16'h5555;
    defparam add_19120_22.INIT1 = 16'h5555;
    defparam add_19120_22.INJECT1_0 = "NO";
    defparam add_19120_22.INJECT1_1 = "NO";
    CCU2D add_19120_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26240), .COUT(n26241));
    defparam add_19120_20.INIT0 = 16'h5555;
    defparam add_19120_20.INIT1 = 16'h5555;
    defparam add_19120_20.INJECT1_0 = "NO";
    defparam add_19120_20.INJECT1_1 = "NO";
    CCU2D add_19120_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26239), .COUT(n26240));
    defparam add_19120_18.INIT0 = 16'h5555;
    defparam add_19120_18.INIT1 = 16'h5555;
    defparam add_19120_18.INJECT1_0 = "NO";
    defparam add_19120_18.INJECT1_1 = "NO";
    CCU2D add_19120_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26238), .COUT(n26239));
    defparam add_19120_16.INIT0 = 16'h5555;
    defparam add_19120_16.INIT1 = 16'h5555;
    defparam add_19120_16.INJECT1_0 = "NO";
    defparam add_19120_16.INJECT1_1 = "NO";
    CCU2D add_19120_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26237), .COUT(n26238));
    defparam add_19120_14.INIT0 = 16'h5555;
    defparam add_19120_14.INIT1 = 16'h5555;
    defparam add_19120_14.INJECT1_0 = "NO";
    defparam add_19120_14.INJECT1_1 = "NO";
    CCU2D add_19120_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26236), .COUT(n26237));
    defparam add_19120_12.INIT0 = 16'h5555;
    defparam add_19120_12.INIT1 = 16'h5555;
    defparam add_19120_12.INJECT1_0 = "NO";
    defparam add_19120_12.INJECT1_1 = "NO";
    CCU2D add_19120_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26235), .COUT(n26236));
    defparam add_19120_10.INIT0 = 16'h5555;
    defparam add_19120_10.INIT1 = 16'h5555;
    defparam add_19120_10.INJECT1_0 = "NO";
    defparam add_19120_10.INJECT1_1 = "NO";
    CCU2D add_19120_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26234), 
          .COUT(n26235));
    defparam add_19120_8.INIT0 = 16'h5555;
    defparam add_19120_8.INIT1 = 16'h5555;
    defparam add_19120_8.INJECT1_0 = "NO";
    defparam add_19120_8.INJECT1_1 = "NO";
    CCU2D add_19120_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26233), 
          .COUT(n26234));
    defparam add_19120_6.INIT0 = 16'h5555;
    defparam add_19120_6.INIT1 = 16'h5555;
    defparam add_19120_6.INJECT1_0 = "NO";
    defparam add_19120_6.INJECT1_1 = "NO";
    CCU2D add_19120_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26232), 
          .COUT(n26233));
    defparam add_19120_4.INIT0 = 16'h5555;
    defparam add_19120_4.INIT1 = 16'h5aaa;
    defparam add_19120_4.INJECT1_0 = "NO";
    defparam add_19120_4.INJECT1_1 = "NO";
    CCU2D add_19120_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26232));
    defparam add_19120_2.INIT0 = 16'h7000;
    defparam add_19120_2.INIT1 = 16'h5aaa;
    defparam add_19120_2.INJECT1_0 = "NO";
    defparam add_19120_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (read_value, \read_value[7]_adj_7 , n46, n3, databus, 
            \read_value[13]_adj_8 , read_value_adj_215, n47, \read_value[7]_adj_41 , 
            n30372, \read_value[13]_adj_42 , n6, databus_out, n32379, 
            n8, \register_addr[0] , \register_addr[1] , n3_adj_43, \select[7] , 
            n30395, n176, n2, \read_value[5]_adj_44 , n3_adj_45, \read_value[11]_adj_46 , 
            \read_value[11]_adj_47 , n6_adj_48, \read_value[11]_adj_49 , 
            n30367, \read_value[26]_adj_50 , read_size, \select[1] , 
            n30454, \reg_size[2] , \sendcount[3] , n4, n3_adj_51, 
            \read_value[13]_adj_52 , \read_value[31]_adj_53 , \register_addr[4] , 
            n30427, \register_addr[5] , n30371, \read_value[31]_adj_54 , 
            n6_adj_55, rw, \read_value[31]_adj_56 , \read_value[6]_adj_57 , 
            n5, prev_select, n32377, n30338, n30374, prev_select_adj_58, 
            n30331, n3_adj_59, \read_value[10]_adj_60 , \read_value[10]_adj_61 , 
            n6_adj_62, n3_adj_63, \read_value[30]_adj_64 , \read_value[30]_adj_65 , 
            n6_adj_66, \read_value[30]_adj_67 , n3_adj_68, \read_value[29]_adj_69 , 
            \read_value[29]_adj_70 , n6_adj_71, \read_value[10]_adj_72 , 
            \read_value[29]_adj_73 , n3_adj_74, \read_value[28]_adj_75 , 
            \read_value[28]_adj_76 , n6_adj_77, \read_value[28]_adj_78 , 
            n8_adj_79, \read_value[6]_adj_80 , n3_adj_81, \read_value[6]_adj_82 , 
            \read_value[27]_adj_83 , n3_adj_84, \read_value[27]_adj_85 , 
            n6_adj_86, \read_value[27]_adj_87 , \read_value[5]_adj_88 , 
            n5_adj_89, n2_adj_90, \read_value[5]_adj_91 , \read_value[26]_adj_92 , 
            n6_adj_93, \read_value[9]_adj_94 , \read_value[26]_adj_95 , 
            n3_adj_96, \read_value[25]_adj_97 , \read_value[9]_adj_98 , 
            n6_adj_99, \register_addr[2] , \read_value[9]_adj_100 , n2_adj_101, 
            \read_value[7]_adj_102 , n5_adj_103, n8_adj_104, \read_value[25]_adj_105 , 
            n6_adj_106, \read_value[25]_adj_107 , n3_adj_108, n2_adj_109, 
            \read_value[24]_adj_110 , \read_value[24]_adj_111 , n6_adj_112, 
            n2_adj_113, \read_value[24]_adj_114 , \read_value[0]_adj_115 , 
            n5_adj_116, n3_adj_117, \read_value[4]_adj_118 , n5_adj_119, 
            n8_adj_120, \read_value[23]_adj_121 , \read_value[4]_adj_122 , 
            \read_value[23]_adj_123 , n6_adj_124, \read_value[23]_adj_125 , 
            n2_adj_126, n3_adj_127, \read_value[4]_adj_128 , \read_value[22]_adj_129 , 
            \read_value[22]_adj_130 , n6_adj_131, \read_value[22]_adj_132 , 
            n3_adj_133, \read_value[21]_adj_134 , \read_value[21]_adj_135 , 
            n6_adj_136, n8_adj_137, \read_value[21]_adj_138 , n3_adj_139, 
            \read_value[20]_adj_140 , \read_value[20]_adj_141 , n6_adj_142, 
            \read_value[20]_adj_143 , n3_adj_144, \read_value[19]_adj_145 , 
            \read_value[19]_adj_146 , n6_adj_147, \read_value[19]_adj_148 , 
            n3_adj_149, \read_value[18]_adj_150 , \read_value[18]_adj_151 , 
            n6_adj_152, \read_value[18]_adj_153 , n3_adj_154, \read_value[17]_adj_155 , 
            \read_value[17]_adj_156 , n6_adj_157, \read_value[17]_adj_158 , 
            n3_adj_159, \read_value[16]_adj_160 , \read_value[16]_adj_161 , 
            n6_adj_162, \read_value[16]_adj_163 , n3_adj_164, \read_value[15]_adj_165 , 
            \read_value[15]_adj_166 , n6_adj_167, \read_value[15]_adj_168 , 
            n3_adj_169, \read_value[14]_adj_170 , \read_value[14]_adj_171 , 
            n6_adj_172, \read_value[14]_adj_173 , n2_adj_174, \read_value[2]_adj_175 , 
            n5_adj_176, n3_adj_177, \read_value[12]_adj_178 , \read_value[12]_adj_179 , 
            n6_adj_180, \read_value[12]_adj_181 , n8_adj_182, n3_adj_183, 
            \read_value[8]_adj_184 , \read_value[8]_adj_185 , n6_adj_186, 
            \read_value[8]_adj_187 , \read_size[0]_adj_188 , n30361, n11, 
            n30396, \read_size[0]_adj_189 , n16, \read_size[0]_adj_190 , 
            \read_size[0]_adj_191 , n30358, n12, \read_size[0]_adj_192 , 
            \read_size[0]_adj_193 , \read_size[0]_adj_194 , n30391, \select[2] , 
            \read_size[2]_adj_195 , \read_value[0]_adj_196 , \read_size[2]_adj_197 , 
            \read_value[1]_adj_198 , \read_value[2]_adj_199 , n4_adj_200, 
            \read_value[2]_adj_201 , \read_value[0]_adj_202 , \read_value[1]_adj_203 , 
            n30339, n2_adj_204, \read_size[2]_adj_205 , \read_size[2]_adj_206 , 
            \read_size[2]_adj_207 , \read_size[2]_adj_208 , \read_value[3]_adj_209 , 
            n5_adj_210, n8_adj_211, \read_value[3]_adj_212 , \read_value[3]_adj_213 , 
            n1, n5_adj_214, GND_net, n28765, debug_c_c, n30303, 
            rc_ch8_c, n26618, n28910, n13624, rc_ch7_c, n26601, 
            n28859, n28775, n14284, rc_ch4_c, n28857, n14306, n28723, 
            n26592, n28855, rc_ch3_c, n26607, n14307, n28770, n28853, 
            n26604, n14308, rc_ch2_c, n28773, n32380, n28851, n14309, 
            rc_ch1_c, n28725, n26596) /* synthesis syn_module_defined=1 */ ;
    input [31:0]read_value;
    input \read_value[7]_adj_7 ;
    input n46;
    input n3;
    output [31:0]databus;
    input \read_value[13]_adj_8 ;
    input [31:0]read_value_adj_215;
    input n47;
    input \read_value[7]_adj_41 ;
    input n30372;
    input \read_value[13]_adj_42 ;
    input n6;
    input [31:0]databus_out;
    input n32379;
    input n8;
    input \register_addr[0] ;
    input \register_addr[1] ;
    input n3_adj_43;
    input \select[7] ;
    input n30395;
    input n176;
    input n2;
    input \read_value[5]_adj_44 ;
    input n3_adj_45;
    input \read_value[11]_adj_46 ;
    input \read_value[11]_adj_47 ;
    input n6_adj_48;
    input \read_value[11]_adj_49 ;
    input n30367;
    input \read_value[26]_adj_50 ;
    input [2:0]read_size;
    input \select[1] ;
    output n30454;
    output \reg_size[2] ;
    input \sendcount[3] ;
    output n4;
    input n3_adj_51;
    input \read_value[13]_adj_52 ;
    input \read_value[31]_adj_53 ;
    input \register_addr[4] ;
    input n30427;
    input \register_addr[5] ;
    output n30371;
    input \read_value[31]_adj_54 ;
    input n6_adj_55;
    input rw;
    input \read_value[31]_adj_56 ;
    input \read_value[6]_adj_57 ;
    input n5;
    input prev_select;
    input n32377;
    output n30338;
    output n30374;
    input prev_select_adj_58;
    output n30331;
    input n3_adj_59;
    input \read_value[10]_adj_60 ;
    input \read_value[10]_adj_61 ;
    input n6_adj_62;
    input n3_adj_63;
    input \read_value[30]_adj_64 ;
    input \read_value[30]_adj_65 ;
    input n6_adj_66;
    input \read_value[30]_adj_67 ;
    input n3_adj_68;
    input \read_value[29]_adj_69 ;
    input \read_value[29]_adj_70 ;
    input n6_adj_71;
    input \read_value[10]_adj_72 ;
    input \read_value[29]_adj_73 ;
    input n3_adj_74;
    input \read_value[28]_adj_75 ;
    input \read_value[28]_adj_76 ;
    input n6_adj_77;
    input \read_value[28]_adj_78 ;
    input n8_adj_79;
    input \read_value[6]_adj_80 ;
    input n3_adj_81;
    input \read_value[6]_adj_82 ;
    input \read_value[27]_adj_83 ;
    input n3_adj_84;
    input \read_value[27]_adj_85 ;
    input n6_adj_86;
    input \read_value[27]_adj_87 ;
    input \read_value[5]_adj_88 ;
    input n5_adj_89;
    input n2_adj_90;
    input \read_value[5]_adj_91 ;
    input \read_value[26]_adj_92 ;
    input n6_adj_93;
    input \read_value[9]_adj_94 ;
    input \read_value[26]_adj_95 ;
    input n3_adj_96;
    input \read_value[25]_adj_97 ;
    input \read_value[9]_adj_98 ;
    input n6_adj_99;
    input \register_addr[2] ;
    input \read_value[9]_adj_100 ;
    input n2_adj_101;
    input \read_value[7]_adj_102 ;
    input n5_adj_103;
    input n8_adj_104;
    input \read_value[25]_adj_105 ;
    input n6_adj_106;
    input \read_value[25]_adj_107 ;
    input n3_adj_108;
    input n2_adj_109;
    input \read_value[24]_adj_110 ;
    input \read_value[24]_adj_111 ;
    input n6_adj_112;
    input n2_adj_113;
    input \read_value[24]_adj_114 ;
    input \read_value[0]_adj_115 ;
    input n5_adj_116;
    input n3_adj_117;
    input \read_value[4]_adj_118 ;
    input n5_adj_119;
    input n8_adj_120;
    input \read_value[23]_adj_121 ;
    input \read_value[4]_adj_122 ;
    input \read_value[23]_adj_123 ;
    input n6_adj_124;
    input \read_value[23]_adj_125 ;
    input n2_adj_126;
    input n3_adj_127;
    input \read_value[4]_adj_128 ;
    input \read_value[22]_adj_129 ;
    input \read_value[22]_adj_130 ;
    input n6_adj_131;
    input \read_value[22]_adj_132 ;
    input n3_adj_133;
    input \read_value[21]_adj_134 ;
    input \read_value[21]_adj_135 ;
    input n6_adj_136;
    input n8_adj_137;
    input \read_value[21]_adj_138 ;
    input n3_adj_139;
    input \read_value[20]_adj_140 ;
    input \read_value[20]_adj_141 ;
    input n6_adj_142;
    input \read_value[20]_adj_143 ;
    input n3_adj_144;
    input \read_value[19]_adj_145 ;
    input \read_value[19]_adj_146 ;
    input n6_adj_147;
    input \read_value[19]_adj_148 ;
    input n3_adj_149;
    input \read_value[18]_adj_150 ;
    input \read_value[18]_adj_151 ;
    input n6_adj_152;
    input \read_value[18]_adj_153 ;
    input n3_adj_154;
    input \read_value[17]_adj_155 ;
    input \read_value[17]_adj_156 ;
    input n6_adj_157;
    input \read_value[17]_adj_158 ;
    input n3_adj_159;
    input \read_value[16]_adj_160 ;
    input \read_value[16]_adj_161 ;
    input n6_adj_162;
    input \read_value[16]_adj_163 ;
    input n3_adj_164;
    input \read_value[15]_adj_165 ;
    input \read_value[15]_adj_166 ;
    input n6_adj_167;
    input \read_value[15]_adj_168 ;
    input n3_adj_169;
    input \read_value[14]_adj_170 ;
    input \read_value[14]_adj_171 ;
    input n6_adj_172;
    input \read_value[14]_adj_173 ;
    input n2_adj_174;
    input \read_value[2]_adj_175 ;
    input n5_adj_176;
    input n3_adj_177;
    input \read_value[12]_adj_178 ;
    input \read_value[12]_adj_179 ;
    input n6_adj_180;
    input \read_value[12]_adj_181 ;
    input n8_adj_182;
    input n3_adj_183;
    input \read_value[8]_adj_184 ;
    input \read_value[8]_adj_185 ;
    input n6_adj_186;
    input \read_value[8]_adj_187 ;
    input \read_size[0]_adj_188 ;
    input n30361;
    output n11;
    input n30396;
    input \read_size[0]_adj_189 ;
    output n16;
    input \read_size[0]_adj_190 ;
    input \read_size[0]_adj_191 ;
    input n30358;
    output n12;
    input \read_size[0]_adj_192 ;
    input \read_size[0]_adj_193 ;
    input \read_size[0]_adj_194 ;
    input n30391;
    input \select[2] ;
    input \read_size[2]_adj_195 ;
    input \read_value[0]_adj_196 ;
    input \read_size[2]_adj_197 ;
    input \read_value[1]_adj_198 ;
    input \read_value[2]_adj_199 ;
    input n4_adj_200;
    input \read_value[2]_adj_201 ;
    input \read_value[0]_adj_202 ;
    input \read_value[1]_adj_203 ;
    input n30339;
    input n2_adj_204;
    input \read_size[2]_adj_205 ;
    input \read_size[2]_adj_206 ;
    input \read_size[2]_adj_207 ;
    input \read_size[2]_adj_208 ;
    input \read_value[3]_adj_209 ;
    input n5_adj_210;
    input n8_adj_211;
    input \read_value[3]_adj_212 ;
    input \read_value[3]_adj_213 ;
    input n1;
    input n5_adj_214;
    input GND_net;
    output n28765;
    input debug_c_c;
    input n30303;
    input rc_ch8_c;
    input n26618;
    output n28910;
    input n13624;
    input rc_ch7_c;
    input n26601;
    output n28859;
    output n28775;
    input n14284;
    input rc_ch4_c;
    output n28857;
    input n14306;
    output n28723;
    input n26592;
    output n28855;
    input rc_ch3_c;
    input n26607;
    input n14307;
    output n28770;
    output n28853;
    input n26604;
    input n14308;
    input rc_ch2_c;
    output n28773;
    input n32380;
    output n28851;
    input n14309;
    input rc_ch1_c;
    output n28725;
    input n26596;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30343, n14, n9, n14_adj_55, n5_c, n30345;
    wire [7:0]read_value_adj_407;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(210[12:22])
    
    wire n46_adj_59, n12_c, n12_adj_61, n6_adj_62_c, n12_adj_63, n16_c;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n30192, n29684, n29683, n29685, n9_adj_64, n14_adj_65, 
        n5_adj_67, n29807, n29314, n30235, n30274, n30198, n29418, 
        n29780;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(211[12:21])
    
    wire n17, n6_adj_69, n16_adj_70;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n29775, n29309, n29774, n14_adj_73, n9_adj_74, n14_adj_75, 
        n5_adj_77, n1016;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n29416, n12_adj_80, n30193;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n29415, n29777, n1001, n29778, n29802, n29801, n29804, 
        n1046, n29805, n30195, n1031, n30196, n9_adj_85, n14_adj_86, 
        n5_adj_88, n30230, n29417, n12_adj_93, n29311, n14_adj_98, 
        n30229, n30232, n30233, n9_adj_101, n14_adj_102, n5_adj_104, 
        n12_adj_107, n9_adj_109, n14_adj_110, n5_adj_112, n12_adj_115, 
        n9_adj_119, n14_adj_120, n5_adj_122, n30269, n12_adj_125, 
        n30268, n9_adj_131, n14_adj_132, n5_adj_134, n12_adj_137, 
        n30271, n986, n30272, n12_adj_142, n9_adj_146, n14_adj_147, 
        n5_adj_149, n9_adj_152, n14_adj_153, n5_adj_155, n12_adj_157, 
        n17_adj_163, n12_adj_167, n29312, n29686, n9_adj_172, n14_adj_173, 
        n5_adj_175, n12_adj_178, n29313, n29310, n17_adj_182, n6_adj_183, 
        n16_adj_184, n12_adj_191, n9_adj_195, n14_adj_196, n5_adj_198, 
        n17_adj_199, n6_adj_200, n16_adj_201, n12_adj_205, n29412, 
        n17_adj_207, n6_adj_208, n16_adj_209, n14_adj_214, n9_adj_216, 
        n14_adj_217, n5_adj_219, n30273, n30270, n14_adj_221, n12_adj_224, 
        n12_adj_230, n16_adj_235, n18, n9_adj_237, n14_adj_238, n5_adj_240, 
        n12_adj_244, n1061, n29687, n9_adj_248, n14_adj_249, n5_adj_251, 
        n12_adj_254, n12_adj_257, n30234, n30231, n9_adj_261, n14_adj_262, 
        n5_adj_264, n30197, n30194, n12_adj_267, n9_adj_271, n14_adj_272, 
        n5_adj_274, n12_adj_277, n9_adj_281, n14_adj_282, n5_adj_284, 
        n12_adj_287, n29413, n9_adj_291, n14_adj_292, n5_adj_294, 
        n12_adj_297, n9_adj_301, n14_adj_302, n5_adj_304, n12_adj_307, 
        n9_adj_311, n14_adj_312, n5_adj_314, n12_adj_317, n9_adj_321, 
        n14_adj_322, n5_adj_324, n12_adj_327, n17_adj_331, n6_adj_332, 
        n16_adj_333, n14_adj_336, n9_adj_338, n14_adj_339, n5_adj_341, 
        n12_adj_344, n12_adj_349, n9_adj_351, n14_adj_352, n5_adj_354, 
        n29308, n12_adj_357, n13, n10, n6_adj_371, n1_c, n21, 
        n14_adj_377, n29689, n11_adj_381, n17_adj_386, n6_adj_387, 
        n16_adj_388, n15, n18_adj_394, n14_adj_396, n12_adj_399, n29806, 
        n29803, n29414, n29779, n29776, n29688;
    
    LUT4 i4_4_lut (.A(read_value[7]), .B(\read_value[7]_adj_7 ), .C(n46), 
         .D(n30343), .Z(n14)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut.init = 16'heca0;
    LUT4 i7_4_lut (.A(n9), .B(n14_adj_55), .C(n3), .D(n5_c), .Z(databus[13])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(\read_value[13]_adj_8 ), .B(read_value_adj_215[13]), 
         .C(n30345), .D(n47), .Z(n9)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i2_4_lut (.A(\read_value[7]_adj_41 ), .B(read_value_adj_407[7]), 
         .C(n30372), .D(n46_adj_59), .Z(n12_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 i6_4_lut (.A(\read_value[13]_adj_42 ), .B(n12_adj_61), .C(n6), 
         .D(n30372), .Z(n14_adj_55)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 Select_4222_i6_2_lut (.A(databus_out[5]), .B(n32379), .Z(n6_adj_62_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4222_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_66 (.A(read_value_adj_215[5]), .B(n12_adj_63), .C(n8), 
         .D(n47), .Z(n16_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_66.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_22277 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n30192)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22277.init = 16'h2222;
    LUT4 Select_4204_i5_2_lut (.A(databus_out[13]), .B(n32379), .Z(n5_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4204_i5_2_lut.init = 16'h2222;
    PFUMX i22068 (.BLUT(n29684), .ALUT(n29683), .C0(\register_addr[1] ), 
          .Z(n29685));
    LUT4 i7_4_lut_adj_67 (.A(n9_adj_64), .B(n14_adj_65), .C(n3_adj_43), 
         .D(n5_adj_67), .Z(databus[26])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_67.init = 16'hfffe;
    FD1S3IX read_value__i6 (.D(n29807), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n29314), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n30235), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i0 (.D(n30274), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n30198), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n29418), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i1 (.D(n29780), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 i9_4_lut (.A(n17), .B(n6_adj_69), .C(n16_adj_70), .D(n2), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 register_addr_1__bdd_2_lut_22084 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n29683)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22084.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_22085 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n29684)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22085.init = 16'he4e4;
    LUT4 register_addr_1__bdd_3_lut_22108 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n29775)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22108.init = 16'he4e4;
    LUT4 register_addr_1__bdd_3_lut_21980 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n29309)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21980.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_22107 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n29774)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22107.init = 16'h2222;
    LUT4 i4_4_lut_adj_68 (.A(read_value[5]), .B(\read_value[5]_adj_44 ), 
         .C(n46), .D(n30343), .Z(n14_adj_73)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_68.init = 16'heca0;
    LUT4 i7_4_lut_adj_69 (.A(n9_adj_74), .B(n14_adj_75), .C(n3_adj_45), 
         .D(n5_adj_77), .Z(databus[11])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_69.init = 16'hfffe;
    LUT4 n1016_bdd_3_lut_22299 (.A(n1016), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n29416)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1016_bdd_3_lut_22299.init = 16'he2e2;
    LUT4 i1_4_lut_adj_70 (.A(\read_value[11]_adj_46 ), .B(read_value_adj_215[11]), 
         .C(n30345), .D(n47), .Z(n9_adj_74)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_70.init = 16'heca0;
    LUT4 i6_4_lut_adj_71 (.A(\read_value[11]_adj_47 ), .B(n12_adj_80), .C(n6_adj_48), 
         .D(n30372), .Z(n14_adj_75)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_71.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_22278 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n30193)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22278.init = 16'he4e4;
    LUT4 Select_4210_i5_2_lut (.A(databus_out[11]), .B(n32379), .Z(n5_adj_77)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4210_i5_2_lut.init = 16'h2222;
    LUT4 n1016_bdd_3_lut_21983 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n29415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1016_bdd_3_lut_21983.init = 16'hcaca;
    LUT4 i4_4_lut_adj_72 (.A(\read_value[11]_adj_49 ), .B(read_value[11]), 
         .C(n30367), .D(n46), .Z(n12_adj_80)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_72.init = 16'heca0;
    LUT4 n1001_bdd_3_lut_22096 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n29777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1001_bdd_3_lut_22096.init = 16'hcaca;
    LUT4 n1001_bdd_3_lut_22305 (.A(n1001), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n29778)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1001_bdd_3_lut_22305.init = 16'he2e2;
    LUT4 register_addr_1__bdd_3_lut_22260 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n29802)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22260.init = 16'he4e4;
    LUT4 i1_4_lut_adj_73 (.A(\read_value[26]_adj_50 ), .B(read_value_adj_215[26]), 
         .C(n30345), .D(n47), .Z(n9_adj_64)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_73.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22259 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n29801)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22259.init = 16'h2222;
    LUT4 n1046_bdd_3_lut_22113 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n29804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1046_bdd_3_lut_22113.init = 16'hcaca;
    LUT4 n1046_bdd_3_lut_22289 (.A(n1046), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n29805)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1046_bdd_3_lut_22289.init = 16'he2e2;
    LUT4 n1031_bdd_3_lut_22265 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n30195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1031_bdd_3_lut_22265.init = 16'hcaca;
    LUT4 n1031_bdd_3_lut_22724 (.A(n1031), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n30196)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1031_bdd_3_lut_22724.init = 16'he2e2;
    LUT4 Select_4236_i1_2_lut_rep_445 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n30454)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4236_i1_2_lut_rep_445.init = 16'h8888;
    LUT4 equal_52_i4_3_lut_4_lut (.A(read_size[1]), .B(\select[1] ), .C(\reg_size[2] ), 
         .D(\sendcount[3] ), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam equal_52_i4_3_lut_4_lut.init = 16'h7f80;
    LUT4 i7_4_lut_adj_74 (.A(n9_adj_85), .B(n14_adj_86), .C(n3_adj_51), 
         .D(n5_adj_88), .Z(databus[31])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_74.init = 16'hfffe;
    LUT4 i4_4_lut_adj_75 (.A(\read_value[13]_adj_52 ), .B(read_value[13]), 
         .C(n30367), .D(n46), .Z(n12_adj_61)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_75.init = 16'heca0;
    LUT4 i1_4_lut_adj_76 (.A(\read_value[31]_adj_53 ), .B(read_value_adj_215[31]), 
         .C(n30345), .D(n47), .Z(n9_adj_85)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_76.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_22294 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n30230)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22294.init = 16'he4e4;
    PFUMX i21984 (.BLUT(n29416), .ALUT(n29415), .C0(\register_addr[1] ), 
          .Z(n29417));
    LUT4 i1_2_lut_rep_362_3_lut (.A(\register_addr[4] ), .B(n30427), .C(\register_addr[5] ), 
         .Z(n30371)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_362_3_lut.init = 16'h8080;
    LUT4 i6_4_lut_adj_77 (.A(\read_value[31]_adj_54 ), .B(n12_adj_93), .C(n6_adj_55), 
         .D(n30372), .Z(n14_adj_86)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_77.init = 16'hfefc;
    LUT4 Select_4150_i5_2_lut (.A(databus_out[31]), .B(rw), .Z(n5_adj_88)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4150_i5_2_lut.init = 16'h2222;
    LUT4 \register_1[[5__bdd_3_lut_22103  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n29311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_22103 .init = 16'hcaca;
    LUT4 i4_4_lut_adj_78 (.A(\read_value[31]_adj_56 ), .B(read_value[31]), 
         .C(n30367), .D(n46), .Z(n12_adj_93)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_78.init = 16'heca0;
    LUT4 i7_4_lut_adj_79 (.A(\read_value[6]_adj_57 ), .B(n14_adj_98), .C(n5), 
         .D(n30345), .Z(n17)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_79.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_22293 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n30229)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22293.init = 16'h2222;
    LUT4 i1_2_lut_rep_329_3_lut_4_lut (.A(\register_addr[4] ), .B(n30427), 
         .C(prev_select), .D(n32377), .Z(n30338)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_329_3_lut_4_lut.init = 16'h0800;
    LUT4 i20_2_lut_rep_336_3_lut_4_lut (.A(\register_addr[4] ), .B(n30427), 
         .C(rw), .D(n32377), .Z(n30345)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20_2_lut_rep_336_3_lut_4_lut.init = 16'h8000;
    LUT4 \register_1[[4__bdd_3_lut_22692  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n30232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_22692 .init = 16'hcaca;
    LUT4 \register_1[[4__bdd_2_lut_22693  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n30233)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_22693 .init = 16'h8888;
    LUT4 i1_2_lut_rep_365_3_lut (.A(\register_addr[4] ), .B(n30427), .C(\register_addr[5] ), 
         .Z(n30374)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_365_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_322_3_lut_4_lut (.A(\register_addr[4] ), .B(n30427), 
         .C(prev_select_adj_58), .D(n32377), .Z(n30331)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_322_3_lut_4_lut.init = 16'h0008;
    LUT4 i20_2_lut_rep_334_3_lut_4_lut (.A(\register_addr[4] ), .B(n30427), 
         .C(n32379), .D(n32377), .Z(n30343)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i20_2_lut_rep_334_3_lut_4_lut.init = 16'h0080;
    LUT4 i7_4_lut_adj_80 (.A(n9_adj_101), .B(n14_adj_102), .C(n3_adj_59), 
         .D(n5_adj_104), .Z(databus[10])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_80.init = 16'hfffe;
    LUT4 i1_4_lut_adj_81 (.A(\read_value[10]_adj_60 ), .B(read_value_adj_215[10]), 
         .C(n30345), .D(n47), .Z(n9_adj_101)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_81.init = 16'heca0;
    LUT4 i6_4_lut_adj_82 (.A(\read_value[10]_adj_61 ), .B(n12_adj_107), 
         .C(n6_adj_62), .D(n30372), .Z(n14_adj_102)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_82.init = 16'hfefc;
    LUT4 Select_4213_i5_2_lut (.A(databus_out[10]), .B(rw), .Z(n5_adj_104)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4213_i5_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_83 (.A(n9_adj_109), .B(n14_adj_110), .C(n3_adj_63), 
         .D(n5_adj_112), .Z(databus[30])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_83.init = 16'hfffe;
    LUT4 i1_4_lut_adj_84 (.A(\read_value[30]_adj_64 ), .B(read_value_adj_215[30]), 
         .C(n30345), .D(n47), .Z(n9_adj_109)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_84.init = 16'heca0;
    LUT4 i6_4_lut_adj_85 (.A(\read_value[30]_adj_65 ), .B(n12_adj_115), 
         .C(n6_adj_66), .D(n30372), .Z(n14_adj_110)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_85.init = 16'hfefc;
    LUT4 Select_4153_i5_2_lut (.A(databus_out[30]), .B(rw), .Z(n5_adj_112)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4153_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_86 (.A(\read_value[30]_adj_67 ), .B(read_value[30]), 
         .C(n30367), .D(n46), .Z(n12_adj_115)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_86.init = 16'heca0;
    LUT4 i7_4_lut_adj_87 (.A(n9_adj_119), .B(n14_adj_120), .C(n3_adj_68), 
         .D(n5_adj_122), .Z(databus[29])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_87.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_22317 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n30269)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22317.init = 16'he4e4;
    LUT4 i1_4_lut_adj_88 (.A(\read_value[29]_adj_69 ), .B(read_value_adj_215[29]), 
         .C(n30345), .D(n47), .Z(n9_adj_119)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_88.init = 16'heca0;
    LUT4 i6_4_lut_adj_89 (.A(\read_value[29]_adj_70 ), .B(n12_adj_125), 
         .C(n6_adj_71), .D(n30372), .Z(n14_adj_120)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_89.init = 16'hfefc;
    LUT4 i4_4_lut_adj_90 (.A(\read_value[10]_adj_72 ), .B(read_value[10]), 
         .C(n30367), .D(n46), .Z(n12_adj_107)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_90.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22316 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n30268)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22316.init = 16'h2222;
    LUT4 Select_4156_i5_2_lut (.A(databus_out[29]), .B(rw), .Z(n5_adj_122)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4156_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_91 (.A(\read_value[29]_adj_73 ), .B(read_value[29]), 
         .C(n30367), .D(n46), .Z(n12_adj_125)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_91.init = 16'heca0;
    LUT4 i7_4_lut_adj_92 (.A(n9_adj_131), .B(n14_adj_132), .C(n3_adj_74), 
         .D(n5_adj_134), .Z(databus[28])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_92.init = 16'hfffe;
    LUT4 i1_4_lut_adj_93 (.A(\read_value[28]_adj_75 ), .B(read_value_adj_215[28]), 
         .C(n30345), .D(n47), .Z(n9_adj_131)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_93.init = 16'heca0;
    LUT4 i6_4_lut_adj_94 (.A(\read_value[28]_adj_76 ), .B(n12_adj_137), 
         .C(n6_adj_77), .D(n30372), .Z(n14_adj_132)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_94.init = 16'hfefc;
    LUT4 Select_4221_i6_2_lut (.A(databus_out[6]), .B(rw), .Z(n6_adj_69)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4221_i6_2_lut.init = 16'h2222;
    LUT4 Select_4159_i5_2_lut (.A(databus_out[28]), .B(rw), .Z(n5_adj_134)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4159_i5_2_lut.init = 16'h2222;
    LUT4 n986_bdd_3_lut_22311 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n30271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n986_bdd_3_lut_22311.init = 16'hcaca;
    LUT4 i4_4_lut_adj_95 (.A(\read_value[28]_adj_78 ), .B(read_value[28]), 
         .C(n30367), .D(n46), .Z(n12_adj_137)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_95.init = 16'heca0;
    LUT4 n986_bdd_3_lut_22643 (.A(n986), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n30272)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n986_bdd_3_lut_22643.init = 16'he2e2;
    LUT4 i6_4_lut_adj_96 (.A(read_value_adj_215[6]), .B(n12_adj_142), .C(n8_adj_79), 
         .D(n47), .Z(n16_adj_70)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_96.init = 16'hfefc;
    LUT4 i4_4_lut_adj_97 (.A(read_value[6]), .B(\read_value[6]_adj_80 ), 
         .C(n46), .D(n30343), .Z(n14_adj_98)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_97.init = 16'heca0;
    LUT4 i7_4_lut_adj_98 (.A(n9_adj_146), .B(n14_adj_147), .C(n3_adj_81), 
         .D(n5_adj_149), .Z(databus[27])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_98.init = 16'hfffe;
    LUT4 i2_4_lut_adj_99 (.A(\read_value[6]_adj_82 ), .B(read_value_adj_407[6]), 
         .C(n30372), .D(n46_adj_59), .Z(n12_adj_142)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_99.init = 16'heca0;
    LUT4 i1_4_lut_adj_100 (.A(\read_value[27]_adj_83 ), .B(read_value_adj_215[27]), 
         .C(n30345), .D(n47), .Z(n9_adj_146)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_100.init = 16'heca0;
    LUT4 i7_4_lut_adj_101 (.A(n9_adj_152), .B(n14_adj_153), .C(n3_adj_84), 
         .D(n5_adj_155), .Z(databus[9])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_101.init = 16'hfffe;
    LUT4 i6_4_lut_adj_102 (.A(\read_value[27]_adj_85 ), .B(n12_adj_157), 
         .C(n6_adj_86), .D(n30372), .Z(n14_adj_147)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_102.init = 16'hfefc;
    LUT4 Select_4162_i5_2_lut (.A(databus_out[27]), .B(rw), .Z(n5_adj_149)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4162_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_103 (.A(\read_value[27]_adj_87 ), .B(read_value[27]), 
         .C(n30367), .D(n46), .Z(n12_adj_157)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_103.init = 16'heca0;
    LUT4 i7_4_lut_adj_104 (.A(\read_value[5]_adj_88 ), .B(n14_adj_73), .C(n5_adj_89), 
         .D(n30345), .Z(n17_adj_163)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_104.init = 16'hfefc;
    LUT4 i9_4_lut_adj_105 (.A(n17_adj_163), .B(n6_adj_62_c), .C(n16_c), 
         .D(n2_adj_90), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_105.init = 16'hfffe;
    LUT4 i2_4_lut_adj_106 (.A(\read_value[5]_adj_91 ), .B(read_value_adj_407[5]), 
         .C(n30372), .D(n46_adj_59), .Z(n12_adj_63)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_106.init = 16'heca0;
    LUT4 i6_4_lut_adj_107 (.A(\read_value[26]_adj_92 ), .B(n12_adj_167), 
         .C(n6_adj_93), .D(n30372), .Z(n14_adj_65)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_107.init = 16'hfefc;
    LUT4 \register_1[[5__bdd_2_lut_22104  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n29312)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_22104 .init = 16'h8888;
    LUT4 i1_4_lut_adj_108 (.A(\read_value[9]_adj_94 ), .B(read_value_adj_215[9]), 
         .C(n30345), .D(n47), .Z(n9_adj_152)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_108.init = 16'heca0;
    LUT4 n1061_bdd_3_lut_22070 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n29686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1061_bdd_3_lut_22070.init = 16'hcaca;
    LUT4 Select_4165_i5_2_lut (.A(databus_out[26]), .B(rw), .Z(n5_adj_67)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4165_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_109 (.A(\read_value[26]_adj_95 ), .B(read_value[26]), 
         .C(n30367), .D(n46), .Z(n12_adj_167)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_109.init = 16'heca0;
    LUT4 i14_2_lut (.A(\select[7] ), .B(rw), .Z(n46_adj_59)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam i14_2_lut.init = 16'h8888;
    LUT4 i7_4_lut_adj_110 (.A(n9_adj_172), .B(n14_adj_173), .C(n3_adj_96), 
         .D(n5_adj_175), .Z(databus[25])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_110.init = 16'hfffe;
    LUT4 i1_4_lut_adj_111 (.A(\read_value[25]_adj_97 ), .B(read_value_adj_215[25]), 
         .C(n30345), .D(n47), .Z(n9_adj_172)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_111.init = 16'heca0;
    LUT4 i6_4_lut_adj_112 (.A(\read_value[9]_adj_98 ), .B(n12_adj_178), 
         .C(n6_adj_99), .D(n30372), .Z(n14_adj_153)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_112.init = 16'hfefc;
    LUT4 Select_4216_i5_2_lut (.A(databus_out[9]), .B(rw), .Z(n5_adj_155)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4216_i5_2_lut.init = 16'h2222;
    L6MUX21 i21956 (.D0(n29313), .D1(n29310), .SD(\register_addr[2] ), 
            .Z(n29314));
    LUT4 i4_4_lut_adj_113 (.A(\read_value[9]_adj_100 ), .B(read_value[9]), 
         .C(n30367), .D(n46), .Z(n12_adj_178)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_113.init = 16'heca0;
    LUT4 i9_4_lut_adj_114 (.A(n17_adj_182), .B(n6_adj_183), .C(n16_adj_184), 
         .D(n2_adj_101), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_114.init = 16'hfffe;
    LUT4 i7_4_lut_adj_115 (.A(\read_value[7]_adj_102 ), .B(n14), .C(n5_adj_103), 
         .D(n30345), .Z(n17_adj_182)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_115.init = 16'hfefc;
    LUT4 Select_4220_i6_2_lut (.A(databus_out[7]), .B(rw), .Z(n6_adj_183)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4220_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_116 (.A(read_value_adj_215[7]), .B(n12_c), .C(n8_adj_104), 
         .D(n47), .Z(n16_adj_184)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_116.init = 16'hfefc;
    LUT4 i6_4_lut_adj_117 (.A(\read_value[25]_adj_105 ), .B(n12_adj_191), 
         .C(n6_adj_106), .D(n30372), .Z(n14_adj_173)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_117.init = 16'hfefc;
    LUT4 Select_4168_i5_2_lut (.A(databus_out[25]), .B(n32379), .Z(n5_adj_175)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4168_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_118 (.A(\read_value[25]_adj_107 ), .B(read_value[25]), 
         .C(n30367), .D(n46), .Z(n12_adj_191)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_118.init = 16'heca0;
    LUT4 i7_4_lut_adj_119 (.A(n9_adj_195), .B(n14_adj_196), .C(n3_adj_108), 
         .D(n5_adj_198), .Z(databus[24])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_119.init = 16'hfffe;
    LUT4 i9_4_lut_adj_120 (.A(n17_adj_199), .B(n6_adj_200), .C(n16_adj_201), 
         .D(n2_adj_109), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_120.init = 16'hfffe;
    LUT4 i1_4_lut_adj_121 (.A(\read_value[24]_adj_110 ), .B(read_value_adj_215[24]), 
         .C(n30345), .D(n47), .Z(n9_adj_195)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_121.init = 16'heca0;
    LUT4 i6_4_lut_adj_122 (.A(\read_value[24]_adj_111 ), .B(n12_adj_205), 
         .C(n6_adj_112), .D(n30372), .Z(n14_adj_196)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_122.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_22064 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n29412)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22064.init = 16'h2222;
    LUT4 i9_4_lut_adj_123 (.A(n17_adj_207), .B(n6_adj_208), .C(n16_adj_209), 
         .D(n2_adj_113), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_123.init = 16'hfffe;
    LUT4 Select_4171_i5_2_lut (.A(databus_out[24]), .B(n32379), .Z(n5_adj_198)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4171_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_124 (.A(\read_value[24]_adj_114 ), .B(read_value[24]), 
         .C(n30367), .D(n46), .Z(n12_adj_205)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_124.init = 16'heca0;
    LUT4 i7_4_lut_adj_125 (.A(\read_value[0]_adj_115 ), .B(n14_adj_214), 
         .C(n5_adj_116), .D(n30345), .Z(n17_adj_207)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_125.init = 16'hfefc;
    LUT4 Select_4227_i6_2_lut (.A(databus_out[0]), .B(rw), .Z(n6_adj_208)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4227_i6_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_126 (.A(n9_adj_216), .B(n14_adj_217), .C(n3_adj_117), 
         .D(n5_adj_219), .Z(databus[23])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_126.init = 16'hfffe;
    L6MUX21 i22314 (.D0(n30273), .D1(n30270), .SD(\register_addr[2] ), 
            .Z(n30274));
    LUT4 i7_4_lut_adj_127 (.A(\read_value[4]_adj_118 ), .B(n14_adj_221), 
         .C(n5_adj_119), .D(n30345), .Z(n17_adj_199)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_127.init = 16'hfefc;
    LUT4 Select_4223_i6_2_lut (.A(databus_out[4]), .B(rw), .Z(n6_adj_200)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4223_i6_2_lut.init = 16'h2222;
    PFUMX i22312 (.BLUT(n30272), .ALUT(n30271), .C0(\register_addr[1] ), 
          .Z(n30273));
    LUT4 i6_4_lut_adj_128 (.A(read_value_adj_215[4]), .B(n12_adj_224), .C(n8_adj_120), 
         .D(n47), .Z(n16_adj_201)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_128.init = 16'hfefc;
    LUT4 i1_4_lut_adj_129 (.A(\read_value[23]_adj_121 ), .B(read_value_adj_215[23]), 
         .C(n30345), .D(n47), .Z(n9_adj_216)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_129.init = 16'heca0;
    LUT4 i4_4_lut_adj_130 (.A(read_value[4]), .B(\read_value[4]_adj_122 ), 
         .C(n46), .D(n30343), .Z(n14_adj_221)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_130.init = 16'heca0;
    LUT4 i6_4_lut_adj_131 (.A(\read_value[23]_adj_123 ), .B(n12_adj_230), 
         .C(n6_adj_124), .D(n30372), .Z(n14_adj_217)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_131.init = 16'hfefc;
    LUT4 Select_4174_i5_2_lut (.A(databus_out[23]), .B(n32379), .Z(n5_adj_219)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4174_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_132 (.A(\read_value[23]_adj_125 ), .B(read_value[23]), 
         .C(n30367), .D(n46), .Z(n12_adj_230)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_132.init = 16'heca0;
    LUT4 i8_4_lut (.A(read_value[1]), .B(n16_adj_235), .C(n2_adj_126), 
         .D(n46), .Z(n18)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut.init = 16'hfefc;
    LUT4 i7_4_lut_adj_133 (.A(n9_adj_237), .B(n14_adj_238), .C(n3_adj_127), 
         .D(n5_adj_240), .Z(databus[22])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_133.init = 16'hfffe;
    LUT4 i2_4_lut_adj_134 (.A(\read_value[4]_adj_128 ), .B(read_value_adj_407[4]), 
         .C(n30372), .D(n46_adj_59), .Z(n12_adj_224)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_134.init = 16'heca0;
    LUT4 i1_4_lut_adj_135 (.A(\read_value[22]_adj_129 ), .B(read_value_adj_215[22]), 
         .C(n30345), .D(n47), .Z(n9_adj_237)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_135.init = 16'heca0;
    LUT4 i6_4_lut_adj_136 (.A(\read_value[22]_adj_130 ), .B(n12_adj_244), 
         .C(n6_adj_131), .D(n30372), .Z(n14_adj_238)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_136.init = 16'hfefc;
    LUT4 Select_4177_i5_2_lut (.A(databus_out[22]), .B(rw), .Z(n5_adj_240)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4177_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_137 (.A(\read_value[22]_adj_132 ), .B(read_value[22]), 
         .C(n30367), .D(n46), .Z(n12_adj_244)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_137.init = 16'heca0;
    LUT4 n1061_bdd_3_lut_22322 (.A(n1061), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n29687)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1061_bdd_3_lut_22322.init = 16'he2e2;
    PFUMX i22309 (.BLUT(n30269), .ALUT(n30268), .C0(\register_addr[1] ), 
          .Z(n30270));
    LUT4 i7_4_lut_adj_138 (.A(n9_adj_248), .B(n14_adj_249), .C(n3_adj_133), 
         .D(n5_adj_251), .Z(databus[21])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_138.init = 16'hfffe;
    LUT4 i1_4_lut_adj_139 (.A(\read_value[21]_adj_134 ), .B(read_value_adj_215[21]), 
         .C(n30345), .D(n47), .Z(n9_adj_248)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_139.init = 16'heca0;
    LUT4 i6_4_lut_adj_140 (.A(\read_value[21]_adj_135 ), .B(n12_adj_254), 
         .C(n6_adj_136), .D(n30372), .Z(n14_adj_249)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_140.init = 16'hfefc;
    LUT4 Select_4180_i5_2_lut (.A(databus_out[21]), .B(n32379), .Z(n5_adj_251)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4180_i5_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_141 (.A(read_value_adj_215[0]), .B(n12_adj_257), .C(n8_adj_137), 
         .D(n47), .Z(n16_adj_209)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_141.init = 16'hfefc;
    LUT4 i4_4_lut_adj_142 (.A(\read_value[21]_adj_138 ), .B(read_value[21]), 
         .C(n30367), .D(n46), .Z(n12_adj_254)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_142.init = 16'heca0;
    L6MUX21 i22285 (.D0(n30234), .D1(n30231), .SD(\register_addr[2] ), 
            .Z(n30235));
    PFUMX i22283 (.BLUT(n30233), .ALUT(n30232), .C0(\register_addr[1] ), 
          .Z(n30234));
    PFUMX i22281 (.BLUT(n30230), .ALUT(n30229), .C0(\register_addr[1] ), 
          .Z(n30231));
    LUT4 i7_4_lut_adj_143 (.A(n9_adj_261), .B(n14_adj_262), .C(n3_adj_139), 
         .D(n5_adj_264), .Z(databus[20])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_143.init = 16'hfffe;
    L6MUX21 i22268 (.D0(n30197), .D1(n30194), .SD(\register_addr[2] ), 
            .Z(n30198));
    LUT4 i1_4_lut_adj_144 (.A(\read_value[20]_adj_140 ), .B(read_value_adj_215[20]), 
         .C(n30345), .D(n47), .Z(n9_adj_261)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_144.init = 16'heca0;
    PFUMX i22266 (.BLUT(n30196), .ALUT(n30195), .C0(\register_addr[1] ), 
          .Z(n30197));
    LUT4 i6_4_lut_adj_145 (.A(\read_value[20]_adj_141 ), .B(n12_adj_267), 
         .C(n6_adj_142), .D(n30372), .Z(n14_adj_262)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_145.init = 16'hfefc;
    LUT4 Select_4183_i5_2_lut (.A(databus_out[20]), .B(n32379), .Z(n5_adj_264)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4183_i5_2_lut.init = 16'h2222;
    PFUMX i22263 (.BLUT(n30193), .ALUT(n30192), .C0(\register_addr[1] ), 
          .Z(n30194));
    LUT4 i4_4_lut_adj_146 (.A(\read_value[20]_adj_143 ), .B(read_value[20]), 
         .C(n30367), .D(n46), .Z(n12_adj_267)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_146.init = 16'heca0;
    LUT4 i7_4_lut_adj_147 (.A(n9_adj_271), .B(n14_adj_272), .C(n3_adj_144), 
         .D(n5_adj_274), .Z(databus[19])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_147.init = 16'hfffe;
    LUT4 i1_4_lut_adj_148 (.A(\read_value[19]_adj_145 ), .B(read_value_adj_215[19]), 
         .C(n30345), .D(n47), .Z(n9_adj_271)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_148.init = 16'heca0;
    LUT4 i6_4_lut_adj_149 (.A(\read_value[19]_adj_146 ), .B(n12_adj_277), 
         .C(n6_adj_147), .D(n30372), .Z(n14_adj_272)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_149.init = 16'hfefc;
    LUT4 Select_4186_i5_2_lut (.A(databus_out[19]), .B(n32379), .Z(n5_adj_274)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4186_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_150 (.A(\read_value[19]_adj_148 ), .B(read_value[19]), 
         .C(n30367), .D(n46), .Z(n12_adj_277)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_150.init = 16'heca0;
    LUT4 i7_4_lut_adj_151 (.A(n9_adj_281), .B(n14_adj_282), .C(n3_adj_149), 
         .D(n5_adj_284), .Z(databus[18])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_151.init = 16'hfffe;
    LUT4 i1_4_lut_adj_152 (.A(\read_value[18]_adj_150 ), .B(read_value_adj_215[18]), 
         .C(n30345), .D(n47), .Z(n9_adj_281)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_152.init = 16'heca0;
    LUT4 i6_4_lut_adj_153 (.A(\read_value[18]_adj_151 ), .B(n12_adj_287), 
         .C(n6_adj_152), .D(n30372), .Z(n14_adj_282)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_153.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_22065 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n29413)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22065.init = 16'he4e4;
    LUT4 Select_4189_i5_2_lut (.A(databus_out[18]), .B(n32379), .Z(n5_adj_284)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4189_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_154 (.A(\read_value[18]_adj_153 ), .B(read_value[18]), 
         .C(n30367), .D(n46), .Z(n12_adj_287)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_154.init = 16'heca0;
    LUT4 i7_4_lut_adj_155 (.A(n9_adj_291), .B(n14_adj_292), .C(n3_adj_154), 
         .D(n5_adj_294), .Z(databus[17])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_155.init = 16'hfffe;
    LUT4 i1_4_lut_adj_156 (.A(\read_value[17]_adj_155 ), .B(read_value_adj_215[17]), 
         .C(n30345), .D(n47), .Z(n9_adj_291)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_156.init = 16'heca0;
    LUT4 i6_4_lut_adj_157 (.A(\read_value[17]_adj_156 ), .B(n12_adj_297), 
         .C(n6_adj_157), .D(n30372), .Z(n14_adj_292)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_157.init = 16'hfefc;
    LUT4 Select_4192_i5_2_lut (.A(databus_out[17]), .B(n32379), .Z(n5_adj_294)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4192_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_158 (.A(\read_value[17]_adj_158 ), .B(read_value[17]), 
         .C(n30367), .D(n46), .Z(n12_adj_297)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_158.init = 16'heca0;
    LUT4 i7_4_lut_adj_159 (.A(n9_adj_301), .B(n14_adj_302), .C(n3_adj_159), 
         .D(n5_adj_304), .Z(databus[16])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_159.init = 16'hfffe;
    LUT4 i1_4_lut_adj_160 (.A(\read_value[16]_adj_160 ), .B(read_value_adj_215[16]), 
         .C(n30345), .D(n47), .Z(n9_adj_301)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_160.init = 16'heca0;
    LUT4 i6_4_lut_adj_161 (.A(\read_value[16]_adj_161 ), .B(n12_adj_307), 
         .C(n6_adj_162), .D(n30372), .Z(n14_adj_302)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_161.init = 16'hfefc;
    LUT4 Select_4195_i5_2_lut (.A(databus_out[16]), .B(n32379), .Z(n5_adj_304)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4195_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_162 (.A(\read_value[16]_adj_163 ), .B(read_value[16]), 
         .C(n30367), .D(n46), .Z(n12_adj_307)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_162.init = 16'heca0;
    LUT4 i7_4_lut_adj_163 (.A(n9_adj_311), .B(n14_adj_312), .C(n3_adj_164), 
         .D(n5_adj_314), .Z(databus[15])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_163.init = 16'hfffe;
    LUT4 i1_4_lut_adj_164 (.A(\read_value[15]_adj_165 ), .B(read_value_adj_215[15]), 
         .C(n30345), .D(n47), .Z(n9_adj_311)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_164.init = 16'heca0;
    LUT4 i6_4_lut_adj_165 (.A(\read_value[15]_adj_166 ), .B(n12_adj_317), 
         .C(n6_adj_167), .D(n30372), .Z(n14_adj_312)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_165.init = 16'hfefc;
    LUT4 Select_4198_i5_2_lut (.A(databus_out[15]), .B(n32379), .Z(n5_adj_314)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4198_i5_2_lut.init = 16'h2222;
    PFUMX i21954 (.BLUT(n29312), .ALUT(n29311), .C0(\register_addr[1] ), 
          .Z(n29313));
    LUT4 i4_4_lut_adj_166 (.A(\read_value[15]_adj_168 ), .B(read_value[15]), 
         .C(n30367), .D(n46), .Z(n12_adj_317)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_166.init = 16'heca0;
    LUT4 i7_4_lut_adj_167 (.A(n9_adj_321), .B(n14_adj_322), .C(n3_adj_169), 
         .D(n5_adj_324), .Z(databus[14])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_167.init = 16'hfffe;
    LUT4 i1_4_lut_adj_168 (.A(\read_value[14]_adj_170 ), .B(read_value_adj_215[14]), 
         .C(n30345), .D(n47), .Z(n9_adj_321)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_168.init = 16'heca0;
    LUT4 i6_4_lut_adj_169 (.A(\read_value[14]_adj_171 ), .B(n12_adj_327), 
         .C(n6_adj_172), .D(n30372), .Z(n14_adj_322)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_169.init = 16'hfefc;
    LUT4 Select_4201_i5_2_lut (.A(databus_out[14]), .B(rw), .Z(n5_adj_324)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4201_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_170 (.A(\read_value[14]_adj_173 ), .B(read_value[14]), 
         .C(n30367), .D(n46), .Z(n12_adj_327)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_170.init = 16'heca0;
    LUT4 i9_4_lut_adj_171 (.A(n17_adj_331), .B(n6_adj_332), .C(n16_adj_333), 
         .D(n2_adj_174), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_171.init = 16'hfffe;
    LUT4 i7_4_lut_adj_172 (.A(\read_value[2]_adj_175 ), .B(n14_adj_336), 
         .C(n5_adj_176), .D(n30345), .Z(n17_adj_331)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_172.init = 16'hfefc;
    LUT4 Select_4225_i6_2_lut (.A(databus_out[2]), .B(n32379), .Z(n6_adj_332)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4225_i6_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_173 (.A(n9_adj_338), .B(n14_adj_339), .C(n3_adj_177), 
         .D(n5_adj_341), .Z(databus[12])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_173.init = 16'hfffe;
    LUT4 i1_4_lut_adj_174 (.A(\read_value[12]_adj_178 ), .B(read_value_adj_215[12]), 
         .C(n30345), .D(n47), .Z(n9_adj_338)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_174.init = 16'heca0;
    LUT4 i6_4_lut_adj_175 (.A(\read_value[12]_adj_179 ), .B(n12_adj_344), 
         .C(n6_adj_180), .D(n30372), .Z(n14_adj_339)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_175.init = 16'hfefc;
    LUT4 Select_4207_i5_2_lut (.A(databus_out[12]), .B(rw), .Z(n5_adj_341)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4207_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_176 (.A(\read_value[12]_adj_181 ), .B(read_value[12]), 
         .C(n30367), .D(n46), .Z(n12_adj_344)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_176.init = 16'heca0;
    LUT4 i6_4_lut_adj_177 (.A(read_value_adj_215[2]), .B(n12_adj_349), .C(n8_adj_182), 
         .D(n47), .Z(n16_adj_333)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_177.init = 16'hfefc;
    LUT4 i7_4_lut_adj_178 (.A(n9_adj_351), .B(n14_adj_352), .C(n3_adj_183), 
         .D(n5_adj_354), .Z(databus[8])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_178.init = 16'hfffe;
    LUT4 i1_4_lut_adj_179 (.A(\read_value[8]_adj_184 ), .B(read_value_adj_215[8]), 
         .C(n30345), .D(n47), .Z(n9_adj_351)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_179.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_21979 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n29308)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21979.init = 16'h2222;
    LUT4 i6_4_lut_adj_180 (.A(\read_value[8]_adj_185 ), .B(n12_adj_357), 
         .C(n6_adj_186), .D(n30372), .Z(n14_adj_352)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_180.init = 16'hfefc;
    LUT4 Select_4219_i5_2_lut (.A(databus_out[8]), .B(rw), .Z(n5_adj_354)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4219_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_181 (.A(\read_value[8]_adj_187 ), .B(read_value[8]), 
         .C(n30367), .D(n46), .Z(n12_adj_357)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_181.init = 16'heca0;
    LUT4 i2_4_lut_adj_182 (.A(read_size[0]), .B(\read_size[0]_adj_188 ), 
         .C(\select[1] ), .D(n30361), .Z(n11)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_182.init = 16'heca0;
    LUT4 i7_4_lut_adj_183 (.A(n13), .B(n30396), .C(n10), .D(\read_size[0]_adj_189 ), 
         .Z(n16)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i7_4_lut_adj_183.init = 16'hfefa;
    LUT4 i3_4_lut (.A(\read_size[0]_adj_190 ), .B(\read_size[0]_adj_191 ), 
         .C(n30371), .D(n30358), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 i4_4_lut_adj_184 (.A(read_size_c[0]), .B(\read_size[0]_adj_192 ), 
         .C(\select[7] ), .D(n30374), .Z(n13)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_184.init = 16'heca0;
    LUT4 i1_4_lut_adj_185 (.A(\read_size[0]_adj_193 ), .B(\read_size[0]_adj_194 ), 
         .C(n30391), .D(\select[2] ), .Z(n10)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_185.init = 16'heca0;
    LUT4 i3_4_lut_adj_186 (.A(n30361), .B(n6_adj_371), .C(n1_c), .D(\read_size[2]_adj_195 ), 
         .Z(\reg_size[2] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_186.init = 16'hfefc;
    LUT4 i4_4_lut_adj_187 (.A(read_value[0]), .B(\read_value[0]_adj_196 ), 
         .C(n46), .D(n30343), .Z(n14_adj_214)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_187.init = 16'heca0;
    LUT4 i2_4_lut_adj_188 (.A(\read_size[2]_adj_197 ), .B(n21), .C(n30358), 
         .D(n30427), .Z(n6_adj_371)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_188.init = 16'heca0;
    LUT4 i4_4_lut_adj_189 (.A(read_value_adj_215[1]), .B(\read_value[1]_adj_198 ), 
         .C(n47), .D(n30343), .Z(n14_adj_377)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_189.init = 16'heca0;
    LUT4 Select_4230_i1_2_lut (.A(read_size[2]), .B(\select[1] ), .Z(n1_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4230_i1_2_lut.init = 16'h8888;
    FD1S3IX read_value__i7 (.D(n29689), .CK(\select[7] ), .CD(n30395), 
            .Q(read_value_adj_407[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=673, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 i4_4_lut_adj_190 (.A(read_value[2]), .B(\read_value[2]_adj_199 ), 
         .C(n46), .D(n30343), .Z(n14_adj_336)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_190.init = 16'heca0;
    LUT4 i6_4_lut_adj_191 (.A(n11_adj_381), .B(n4_adj_200), .C(databus_out[1]), 
         .D(rw), .Z(n16_adj_235)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i6_4_lut_adj_191.init = 16'heefe;
    LUT4 i2_4_lut_adj_192 (.A(\read_value[2]_adj_201 ), .B(read_value_adj_407[2]), 
         .C(n30372), .D(n46_adj_59), .Z(n12_adj_349)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_192.init = 16'heca0;
    LUT4 i2_4_lut_adj_193 (.A(\read_value[0]_adj_202 ), .B(read_value_adj_407[0]), 
         .C(n30372), .D(n46_adj_59), .Z(n12_adj_257)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_193.init = 16'heca0;
    LUT4 i1_4_lut_adj_194 (.A(\read_value[1]_adj_203 ), .B(read_value_adj_407[1]), 
         .C(n30339), .D(n46_adj_59), .Z(n11_adj_381)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_194.init = 16'heca0;
    LUT4 i9_4_lut_adj_195 (.A(n17_adj_386), .B(n6_adj_387), .C(n16_adj_388), 
         .D(n2_adj_204), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_195.init = 16'hfffe;
    LUT4 i35_3_lut (.A(\read_size[2]_adj_205 ), .B(\read_size[2]_adj_206 ), 
         .C(\register_addr[4] ), .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i35_3_lut.init = 16'hcaca;
    LUT4 i34_3_lut (.A(\read_size[2]_adj_207 ), .B(\read_size[2]_adj_208 ), 
         .C(\register_addr[4] ), .Z(n18_adj_394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i34_3_lut.init = 16'hcaca;
    LUT4 i7_4_lut_adj_196 (.A(\read_value[3]_adj_209 ), .B(n14_adj_396), 
         .C(n5_adj_210), .D(n30345), .Z(n17_adj_386)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_196.init = 16'hfefc;
    LUT4 Select_4224_i6_2_lut (.A(databus_out[3]), .B(n32379), .Z(n6_adj_387)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4224_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_197 (.A(read_value_adj_215[3]), .B(n12_adj_399), .C(n8_adj_211), 
         .D(n47), .Z(n16_adj_388)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_197.init = 16'hfefc;
    L6MUX21 i22116 (.D0(n29806), .D1(n29803), .SD(\register_addr[2] ), 
            .Z(n29807));
    PFUMX i22114 (.BLUT(n29805), .ALUT(n29804), .C0(\register_addr[1] ), 
          .Z(n29806));
    LUT4 i4_4_lut_adj_198 (.A(read_value[3]), .B(\read_value[3]_adj_212 ), 
         .C(n46), .D(n30343), .Z(n14_adj_396)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_198.init = 16'heca0;
    LUT4 i2_4_lut_adj_199 (.A(\read_value[3]_adj_213 ), .B(read_value_adj_407[3]), 
         .C(n30372), .D(n46_adj_59), .Z(n12_adj_399)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_199.init = 16'heca0;
    LUT4 i9_4_lut_adj_200 (.A(n1), .B(n18), .C(n14_adj_377), .D(n5_adj_214), 
         .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_200.init = 16'hfffe;
    PFUMX i22111 (.BLUT(n29802), .ALUT(n29801), .C0(\register_addr[1] ), 
          .Z(n29803));
    L6MUX21 i21986 (.D0(n29417), .D1(n29414), .SD(\register_addr[2] ), 
            .Z(n29418));
    L6MUX21 i22099 (.D0(n29779), .D1(n29776), .SD(\register_addr[2] ), 
            .Z(n29780));
    PFUMX i22097 (.BLUT(n29778), .ALUT(n29777), .C0(\register_addr[1] ), 
          .Z(n29779));
    PFUMX i22094 (.BLUT(n29775), .ALUT(n29774), .C0(\register_addr[1] ), 
          .Z(n29776));
    PFUMX i36 (.BLUT(n15), .ALUT(n18_adj_394), .C0(\register_addr[5] ), 
          .Z(n21));
    PFUMX i21952 (.BLUT(n29309), .ALUT(n29308), .C0(\register_addr[1] ), 
          .Z(n29310));
    PFUMX i21981 (.BLUT(n29413), .ALUT(n29412), .C0(\register_addr[1] ), 
          .Z(n29414));
    L6MUX21 i22073 (.D0(n29688), .D1(n29685), .SD(\register_addr[2] ), 
            .Z(n29689));
    PFUMX i22071 (.BLUT(n29687), .ALUT(n29686), .C0(\register_addr[1] ), 
          .Z(n29688));
    PWMReceiver recv_ch8 (.GND_net(GND_net), .n28765(n28765), .debug_c_c(debug_c_c), 
            .n30303(n30303), .rc_ch8_c(rc_ch8_c), .n1061(n1061), .n26618(n26618), 
            .n28910(n28910), .\register[6] ({\register[6] }), .n13624(n13624)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(257[14] 261[36])
    PWMReceiver_U1 recv_ch7 (.debug_c_c(debug_c_c), .n30303(n30303), .rc_ch7_c(rc_ch7_c), 
            .GND_net(GND_net), .n1046(n1046), .n26601(n26601), .n28859(n28859), 
            .n28775(n28775), .\register[5] ({\register[5] }), .n14284(n14284)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(252[14] 256[36])
    PWMReceiver_U2 recv_ch4 (.debug_c_c(debug_c_c), .n30303(n30303), .rc_ch4_c(rc_ch4_c), 
            .GND_net(GND_net), .n28857(n28857), .\register[4] ({\register[4] }), 
            .n14306(n14306), .n28723(n28723), .n1031(n1031), .n26592(n26592)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(247[14] 251[36])
    PWMReceiver_U3 recv_ch3 (.n28855(n28855), .n30303(n30303), .debug_c_c(debug_c_c), 
            .rc_ch3_c(rc_ch3_c), .GND_net(GND_net), .n1016(n1016), .n26607(n26607), 
            .\register[3] ({\register[3] }), .n14307(n14307), .n28770(n28770)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(242[14] 246[36])
    PWMReceiver_U4 recv_ch2 (.GND_net(GND_net), .n28853(n28853), .n30303(n30303), 
            .n1001(n1001), .debug_c_c(debug_c_c), .n26604(n26604), .\register[2] ({\register[2] }), 
            .n14308(n14308), .rc_ch2_c(rc_ch2_c), .n28773(n28773)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(237[14] 241[36])
    PWMReceiver_U5 recv_ch1 (.debug_c_c(debug_c_c), .n30303(n30303), .GND_net(GND_net), 
            .n32380(n32380), .n28851(n28851), .\register[1] ({\register[1] }), 
            .n14309(n14309), .rc_ch1_c(rc_ch1_c), .n28725(n28725), .n986(n986), 
            .n26596(n26596)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(232[17] 236[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (GND_net, n28765, debug_c_c, n30303, rc_ch8_c, 
            n1061, n26618, n28910, \register[6] , n13624) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n28765;
    input debug_c_c;
    input n30303;
    input rc_ch8_c;
    output n1061;
    input n26618;
    output n28910;
    output [7:0]\register[6] ;
    input n13624;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25541;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n5;
    wire [15:0]n116;
    
    wire n25542, n26469, n30352, n26804, n30328, n28316, n25540, 
        n25539, n30438, n26768, n26617, n30404, n30439, n30440, 
        n28222, n1067, n1055, n13265, n28317, n30377, n114, n4, 
        n30442, n28423, n30403, n30376, n30443, n30405, n30378, 
        n28529, n28325, n28577, n54, n23, n30353, n28270, n10, 
        n28102, n26665, n6, n28040, n16316, n24;
    wire [7:0]n959;
    wire [7:0]n43;
    
    wire n28209, n25818, n25817, n25816, n25815, n25543, n25546, 
        n25545, n25544;
    
    CCU2D add_1760_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25541), 
          .COUT(n25542), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_7.INIT0 = 16'hd222;
    defparam add_1760_7.INIT1 = 16'hd222;
    defparam add_1760_7.INJECT1_0 = "NO";
    defparam add_1760_7.INJECT1_1 = "NO";
    LUT4 i21791_3_lut_3_lut_4_lut (.A(n26469), .B(n30352), .C(n26804), 
         .D(n30328), .Z(n28316)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i21791_3_lut_3_lut_4_lut.init = 16'h000e;
    CCU2D add_1760_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25540), 
          .COUT(n25541), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_5.INIT0 = 16'hd222;
    defparam add_1760_5.INIT1 = 16'hd222;
    defparam add_1760_5.INJECT1_0 = "NO";
    defparam add_1760_5.INJECT1_1 = "NO";
    CCU2D add_1760_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25539), 
          .COUT(n25540), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_3.INIT0 = 16'hd222;
    defparam add_1760_3.INIT1 = 16'hd222;
    defparam add_1760_3.INJECT1_0 = "NO";
    defparam add_1760_3.INJECT1_1 = "NO";
    LUT4 i21713_4_lut (.A(n30438), .B(n5), .C(n26768), .D(n26617), .Z(n28765)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i21713_4_lut.init = 16'h3233;
    LUT4 i2_3_lut_4_lut (.A(count[0]), .B(n30404), .C(n30439), .D(n30440), 
         .Z(n28222)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n30303), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1067));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_429 (.A(count[15]), .B(count[14]), .Z(n30438)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_429.init = 16'heeee;
    FD1P3AX prev_in_46 (.D(n1067), .SP(n30303), .CK(debug_c_c), .Q(n1055));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(n1055), .B(n1067), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_4_lut_adj_49 (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n13265)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_49.init = 16'hfffe;
    LUT4 i1_2_lut_rep_319_3_lut (.A(count[15]), .B(count[14]), .C(n26768), 
         .Z(n30328)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_319_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n26768), 
         .Z(n28317)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_430 (.A(count[1]), .B(count[2]), .Z(n30439)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_430.init = 16'h8888;
    LUT4 i2_2_lut_rep_368_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(n30440), 
         .D(count[8]), .Z(n30377)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_rep_368_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n114)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_50 (.A(count[1]), .B(count[2]), .C(count[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_50.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_431 (.A(count[6]), .B(count[7]), .Z(n30440)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_431.init = 16'h8888;
    LUT4 i21276_2_lut_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(n30442), 
         .D(count[3]), .Z(n28423)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21276_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_394_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n30403)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_394_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_433 (.A(count[4]), .B(count[5]), .Z(n30442)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_433.init = 16'h8888;
    LUT4 i1_2_lut_rep_395_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n30404)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_395_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_367_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n30376)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_367_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_434 (.A(count[11]), .B(count[10]), .Z(n30443)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_434.init = 16'heeee;
    LUT4 i1_2_lut_rep_396_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n30405)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_396_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_369_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n13265), 
         .D(count[9]), .Z(n30378)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_369_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(n28529), .B(n28325), .C(n30443), .D(n28577), .Z(n26617)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccce;
    LUT4 i21424_4_lut (.A(n54), .B(n13265), .C(n23), .D(n30353), .Z(n28577)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21424_4_lut.init = 16'hfffe;
    FD1P3IX valid_48 (.D(n28316), .SP(n26618), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1061));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_51 (.A(count[8]), .B(n30440), .C(count[0]), 
         .D(n30439), .Z(n28270)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut_adj_51.init = 16'h8000;
    LUT4 i1_2_lut_rep_343_3_lut_4_lut (.A(count[9]), .B(n30443), .C(count[8]), 
         .D(n13265), .Z(n30352)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_343_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_1760_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28317), .B1(n1067), .C1(count[0]), .D1(n1055), .COUT(n25539), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_1.INIT0 = 16'hF000;
    defparam add_1760_1.INIT1 = 16'ha565;
    defparam add_1760_1.INJECT1_0 = "NO";
    defparam add_1760_1.INJECT1_1 = "NO";
    LUT4 i21858_4_lut (.A(n54), .B(n28325), .C(n23), .D(n10), .Z(n28910)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21858_4_lut.init = 16'h3332;
    LUT4 i3_4_lut (.A(count[6]), .B(count[8]), .C(count[7]), .D(n28102), 
         .Z(n26665)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_52 (.A(count[2]), .B(n30442), .C(n6), .D(count[0]), 
         .Z(n28102)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_52.init = 16'hccc8;
    LUT4 i3_4_lut_adj_53 (.A(n30438), .B(n28040), .C(n30443), .D(n30303), 
         .Z(n16316)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_53.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[13]), .B(n24), .C(count[12]), .D(n28325), 
         .Z(n28040)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i2_2_lut (.A(count[3]), .B(count[1]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i31_4_lut (.A(n30376), .B(n26665), .C(count[9]), .D(n30377), 
         .Z(n24)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_4_lut.init = 16'h3a30;
    LUT4 i2_4_lut (.A(n30440), .B(count[5]), .C(count[4]), .D(n4), .Z(n26469)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i21_4_lut (.A(n30404), .B(n26804), .C(n30378), .D(n28270), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_4_lut_adj_54 (.A(count[8]), .B(n30378), .C(n30439), .D(n28423), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_54.init = 16'h0222;
    LUT4 i1_2_lut (.A(n23), .B(n959[7]), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_55 (.A(n23), .B(n959[6]), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_55.init = 16'h8888;
    LUT4 i1_2_lut_adj_56 (.A(n23), .B(n959[5]), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_56.init = 16'h8888;
    LUT4 i1_2_lut_adj_57 (.A(n1067), .B(n1055), .Z(n28325)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_57.init = 16'hbbbb;
    LUT4 i1_2_lut_adj_58 (.A(n23), .B(n959[4]), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_58.init = 16'h8888;
    LUT4 i2_4_lut_adj_59 (.A(count[13]), .B(count[12]), .C(n28209), .D(n30405), 
         .Z(n26768)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_59.init = 16'h8880;
    CCU2D sub_67_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25818), 
          .S0(n959[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_67_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_67_add_2_9.INIT1 = 16'h0000;
    defparam sub_67_add_2_9.INJECT1_0 = "NO";
    defparam sub_67_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_67_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25817), 
          .COUT(n25818), .S0(n959[5]), .S1(n959[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_67_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_67_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_67_add_2_7.INJECT1_0 = "NO";
    defparam sub_67_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_60 (.A(n23), .B(n959[3]), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_60.init = 16'h8888;
    LUT4 i1_2_lut_adj_61 (.A(n23), .B(n959[2]), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_61.init = 16'h8888;
    CCU2D sub_67_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25816), 
          .COUT(n25817), .S0(n959[3]), .S1(n959[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_67_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_67_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_67_add_2_5.INJECT1_0 = "NO";
    defparam sub_67_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_67_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25815), 
          .COUT(n25816), .S0(n959[1]), .S1(n959[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_67_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_67_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_67_add_2_3.INJECT1_0 = "NO";
    defparam sub_67_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_62 (.A(n23), .B(n959[1]), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_62.init = 16'h8888;
    LUT4 i1_4_lut_adj_63 (.A(count[4]), .B(n30403), .C(n114), .D(count[5]), 
         .Z(n28209)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_63.init = 16'hccc8;
    CCU2D sub_67_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25815), 
          .S1(n959[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_67_add_2_1.INIT0 = 16'hF000;
    defparam sub_67_add_2_1.INIT1 = 16'h5555;
    defparam sub_67_add_2_1.INJECT1_0 = "NO";
    defparam sub_67_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_64 (.A(n23), .B(n959[0]), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_64.init = 16'h8888;
    CCU2D add_1760_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25542), 
          .COUT(n25543), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_9.INIT0 = 16'hd222;
    defparam add_1760_9.INIT1 = 16'hd222;
    defparam add_1760_9.INJECT1_0 = "NO";
    defparam add_1760_9.INJECT1_1 = "NO";
    LUT4 i21380_3_lut_4_lut (.A(count[8]), .B(n30378), .C(n26469), .D(n28222), 
         .Z(n28529)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i21380_3_lut_4_lut.init = 16'hfeee;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n30378), .C(n28222), 
         .D(n26469), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i15334_2_lut_rep_344 (.A(count[9]), .B(n26665), .Z(n30353)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i15334_2_lut_rep_344.init = 16'h8888;
    LUT4 i2_3_lut_4_lut_adj_65 (.A(count[9]), .B(n26665), .C(n30443), 
         .D(n13265), .Z(n26804)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_4_lut_adj_65.init = 16'hfff8;
    CCU2D add_1760_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25546), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_17.INIT0 = 16'hd222;
    defparam add_1760_17.INIT1 = 16'h0000;
    defparam add_1760_17.INJECT1_0 = "NO";
    defparam add_1760_17.INJECT1_1 = "NO";
    CCU2D add_1760_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25545), 
          .COUT(n25546), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_15.INIT0 = 16'hd222;
    defparam add_1760_15.INIT1 = 16'hd222;
    defparam add_1760_15.INJECT1_0 = "NO";
    defparam add_1760_15.INJECT1_1 = "NO";
    CCU2D add_1760_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25544), 
          .COUT(n25545), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_13.INIT0 = 16'hd222;
    defparam add_1760_13.INIT1 = 16'hd222;
    defparam add_1760_13.INJECT1_0 = "NO";
    defparam add_1760_13.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13624), .PD(n16316), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1760_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25543), 
          .COUT(n25544), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1760_11.INIT0 = 16'hd222;
    defparam add_1760_11.INIT1 = 16'hd222;
    defparam add_1760_11.INJECT1_0 = "NO";
    defparam add_1760_11.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (debug_c_c, n30303, rc_ch7_c, GND_net, n1046, 
            n26601, n28859, n28775, \register[5] , n14284) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30303;
    input rc_ch7_c;
    input GND_net;
    output n1046;
    input n26601;
    output n28859;
    output n28775;
    output [7:0]\register[5] ;
    input n14284;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n1052, n25552;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n5;
    wire [15:0]n116;
    
    wire n25553, n25551, n28304, n1040, n152, n103, n154, n26373, 
        n30364, n28433, n30337, n13127, n30388, n30387, n30363, 
        n25550, n30461, n30470, n25549, n5_adj_49, n30471, n26769, 
        n28305, n30472, n30415, n30473, n6, n4, n4_adj_50, n54, 
        n28343, n10, n11, n28573, n16259, n28100, n25548, n5_adj_51, 
        n25822;
    wire [7:0]n950;
    
    wire n25821, n25820, n25819;
    wire [7:0]n43;
    
    wire n25547, n26599, n28543, n28361, n4_adj_52, n6_adj_53, n25554;
    
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n30303), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1052));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    CCU2D add_1756_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25552), 
          .COUT(n25553), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_13.INIT0 = 16'hd222;
    defparam add_1756_13.INIT1 = 16'hd222;
    defparam add_1756_13.INJECT1_0 = "NO";
    defparam add_1756_13.INJECT1_1 = "NO";
    CCU2D add_1756_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25551), 
          .COUT(n25552), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_11.INIT0 = 16'hd222;
    defparam add_1756_11.INIT1 = 16'hd222;
    defparam add_1756_11.INJECT1_0 = "NO";
    defparam add_1756_11.INJECT1_1 = "NO";
    FD1P3IX valid_48 (.D(n28304), .SP(n26601), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1046));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1052), .SP(n30303), .CK(debug_c_c), .Q(n1040));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    PFUMX i13749 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    LUT4 i21789_3_lut_3_lut_4_lut (.A(n26373), .B(n30364), .C(n28433), 
         .D(n30337), .Z(n28304)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i21789_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_2_lut_rep_379 (.A(count[9]), .B(n13127), .Z(n30388)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_379.init = 16'heeee;
    LUT4 i1_3_lut_rep_354_4_lut (.A(count[9]), .B(n13127), .C(n30387), 
         .D(count[8]), .Z(n30363)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_3_lut_rep_354_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_355_3_lut (.A(count[9]), .B(n13127), .C(count[8]), 
         .Z(n30364)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_355_3_lut.init = 16'hfefe;
    CCU2D add_1756_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25550), 
          .COUT(n25551), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_9.INIT0 = 16'hd222;
    defparam add_1756_9.INIT1 = 16'hd222;
    defparam add_1756_9.INJECT1_0 = "NO";
    defparam add_1756_9.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_452 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n30461)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_452.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[8]), .D(n30470), 
         .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    CCU2D add_1756_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25549), 
          .COUT(n25550), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_7.INIT0 = 16'hd222;
    defparam add_1756_7.INIT1 = 16'hd222;
    defparam add_1756_7.INJECT1_0 = "NO";
    defparam add_1756_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_461 (.A(count[4]), .B(count[5]), .Z(n30470)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_461.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n5_adj_49)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_462 (.A(count[15]), .B(count[14]), .Z(n30471)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_462.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_42 (.A(count[15]), .B(count[14]), .C(n5), 
         .D(n26769), .Z(n28305)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_42.init = 16'hfffe;
    LUT4 i1_2_lut_rep_328_3_lut (.A(count[15]), .B(count[14]), .C(n26769), 
         .Z(n30337)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_328_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_463 (.A(count[7]), .B(count[6]), .Z(n30472)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_463.init = 16'h8888;
    LUT4 i1_2_lut_rep_406_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n30415)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_406_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n30473), 
         .D(count[8]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_464 (.A(count[2]), .B(count[1]), .Z(n30473)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_464.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4_adj_50)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i21807_4_lut (.A(n54), .B(n28343), .C(n30363), .D(n10), .Z(n28859)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21807_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n30303), .B(n30471), .C(n11), .D(n28573), .Z(n16259)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i4_4_lut (.A(n28100), .B(n28343), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i21420_4_lut (.A(count[12]), .B(count[13]), .C(count[11]), .D(count[10]), 
         .Z(n28573)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21420_4_lut.init = 16'hfffe;
    CCU2D add_1756_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25548), 
          .COUT(n25549), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_5.INIT0 = 16'hd222;
    defparam add_1756_5.INIT1 = 16'hd222;
    defparam add_1756_5.INJECT1_0 = "NO";
    defparam add_1756_5.INJECT1_1 = "NO";
    LUT4 i3_3_lut_rep_378_4_lut (.A(count[3]), .B(n30470), .C(n30472), 
         .D(n30473), .Z(n30387)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_3_lut_rep_378_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(n1040), .B(n1052), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_4_lut_adj_43 (.A(n30388), .B(count[8]), .C(n30387), 
         .D(n54), .Z(n5_adj_51)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_43.init = 16'h00fb;
    CCU2D sub_66_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25822), 
          .S0(n950[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_66_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_66_add_2_9.INIT1 = 16'h0000;
    defparam sub_66_add_2_9.INJECT1_0 = "NO";
    defparam sub_66_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_66_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25821), 
          .COUT(n25822), .S0(n950[5]), .S1(n950[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_66_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_66_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_66_add_2_7.INJECT1_0 = "NO";
    defparam sub_66_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_66_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25820), 
          .COUT(n25821), .S0(n950[3]), .S1(n950[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_66_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_66_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_66_add_2_5.INJECT1_0 = "NO";
    defparam sub_66_add_2_5.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    CCU2D sub_66_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25819), 
          .COUT(n25820), .S0(n950[1]), .S1(n950[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_66_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_66_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_66_add_2_3.INJECT1_0 = "NO";
    defparam sub_66_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_66_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25819), 
          .S1(n950[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_66_add_2_1.INIT0 = 16'hF000;
    defparam sub_66_add_2_1.INIT1 = 16'h5555;
    defparam sub_66_add_2_1.INJECT1_0 = "NO";
    defparam sub_66_add_2_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    LUT4 i15118_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15118_2_lut_4_lut.init = 16'h0400;
    CCU2D add_1756_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25547), 
          .COUT(n25548), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_3.INIT0 = 16'hd222;
    defparam add_1756_3.INIT1 = 16'hd222;
    defparam add_1756_3.INJECT1_0 = "NO";
    defparam add_1756_3.INJECT1_1 = "NO";
    CCU2D add_1756_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28305), .B1(n1052), .C1(count[0]), .D1(n1040), .COUT(n25547), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_1.INIT0 = 16'hF000;
    defparam add_1756_1.INIT1 = 16'ha565;
    defparam add_1756_1.INJECT1_0 = "NO";
    defparam add_1756_1.INJECT1_1 = "NO";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    LUT4 i21723_4_lut (.A(n30471), .B(n5), .C(n26769), .D(n26599), .Z(n28775)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i21723_4_lut.init = 16'h3233;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n5_adj_51), .B(n28343), .C(n28543), .D(n28433), 
         .Z(n26599)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i21286_3_lut (.A(n13127), .B(count[9]), .C(n154), .Z(n28433)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i21286_3_lut.init = 16'heaea;
    LUT4 i3_4_lut (.A(count[12]), .B(n30471), .C(count[13]), .D(n28361), 
         .Z(n13127)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_44 (.A(n30472), .B(count[5]), .C(count[3]), .D(n4), 
         .Z(n26373)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_44.init = 16'h8880;
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n28361)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(n5_adj_49), .B(n28433), .C(n30388), .D(n6), .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_2_lut_adj_45 (.A(n1052), .B(n1040), .Z(n28343)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_45.init = 16'hbbbb;
    LUT4 i2_4_lut_adj_46 (.A(count[13]), .B(count[12]), .C(n28361), .D(n4_adj_52), 
         .Z(n26769)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_46.init = 16'h8880;
    LUT4 i1_4_lut_adj_47 (.A(count[9]), .B(count[4]), .C(n30415), .D(n4_adj_50), 
         .Z(n4_adj_52)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_47.init = 16'hfaea;
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i15117_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15117_2_lut_4_lut.init = 16'h0400;
    LUT4 i23_4_lut (.A(n30461), .B(count[2]), .C(n30470), .D(n6_adj_53), 
         .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i15116_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15116_2_lut_4_lut.init = 16'h0400;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6_adj_53)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i15115_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15115_2_lut_4_lut.init = 16'h0400;
    LUT4 i15114_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15114_2_lut_4_lut.init = 16'h0400;
    LUT4 i15113_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15113_2_lut_4_lut.init = 16'h0400;
    LUT4 i15112_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15112_2_lut_4_lut.init = 16'h0400;
    LUT4 i14877_2_lut_4_lut (.A(n30388), .B(count[8]), .C(n30387), .D(n950[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14877_2_lut_4_lut.init = 16'h0400;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[0]), .B(n30387), .C(n30364), 
         .D(n26373), .Z(n10)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0700;
    LUT4 i21391_3_lut_4_lut (.A(count[0]), .B(n30387), .C(n26373), .D(n30364), 
         .Z(n28543)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21391_3_lut_4_lut.init = 16'hff80;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14284), .PD(n16259), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_48 (.A(count[0]), .B(n30387), .C(count[8]), 
         .Z(n28100)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_48.init = 16'h8080;
    CCU2D add_1756_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25554), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_17.INIT0 = 16'hd222;
    defparam add_1756_17.INIT1 = 16'h0000;
    defparam add_1756_17.INJECT1_0 = "NO";
    defparam add_1756_17.INJECT1_1 = "NO";
    CCU2D add_1756_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25553), 
          .COUT(n25554), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1756_15.INIT0 = 16'hd222;
    defparam add_1756_15.INIT1 = 16'hd222;
    defparam add_1756_15.INJECT1_0 = "NO";
    defparam add_1756_15.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (debug_c_c, n30303, rc_ch4_c, GND_net, n28857, 
            \register[4] , n14306, n28723, n1031, n26592) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30303;
    input rc_ch4_c;
    input GND_net;
    output n28857;
    output [7:0]\register[4] ;
    input n14306;
    output n28723;
    output n1031;
    input n26592;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n20243;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n30459, n30484, n30393, n30392;
    wire [7:0]n941;
    wire [7:0]n43;
    
    wire n13181, n28286, n30332, n1025, n1037, n152, n103, n154, 
        n30458, n30425, n13179, n30368, n30369, n30482, n28377, 
        n30483, n28587, n28146, n30485, n28226, n4, n162, n4_adj_47, 
        n54, n28337, n10, n11, n16272, n26341, n28431;
    wire [15:0]n116;
    
    wire n25826, n25825, n25824, n25823, n25562, n25561, n25560, 
        n25559, n25558, n28021, n28020, n4_adj_48, n28378, n25557, 
        n6, n25556, n25555;
    
    LUT4 i2_2_lut_rep_384_4_lut (.A(n20243), .B(count[3]), .C(n30459), 
         .D(n30484), .Z(n30393)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut_rep_384_4_lut.init = 16'h8000;
    LUT4 i15103_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15103_2_lut_4_lut.init = 16'h0400;
    LUT4 i14871_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14871_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_4_lut_rep_323 (.A(n13181), .B(count[13]), .C(count[12]), .D(n28286), 
         .Z(n30332)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_323.init = 16'heaaa;
    FD1P3AX prev_in_46 (.D(n1037), .SP(n30303), .CK(debug_c_c), .Q(n1025));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n30303), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1037));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    PFUMX i13843 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    LUT4 i2_3_lut_rep_449 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n30458)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_449.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[8]), .D(n30459), 
         .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_450 (.A(count[4]), .B(count[5]), .Z(n30459)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_450.init = 16'h8888;
    LUT4 i1_3_lut_rep_416_4_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .D(n20243), .Z(n30425)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_rep_416_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_383 (.A(count[9]), .B(n13179), .Z(n30392)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_383.init = 16'heeee;
    LUT4 i1_2_lut_rep_359_3_lut (.A(count[9]), .B(n13179), .C(count[8]), 
         .Z(n30368)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_359_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_360_4_lut (.A(count[9]), .B(n13179), .C(n30393), 
         .D(count[8]), .Z(n30369)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i2_3_lut_rep_360_4_lut.init = 16'hfeff;
    LUT4 i5_2_lut_rep_473 (.A(n1025), .B(n1037), .Z(n30482)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_473.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n1025), .B(n1037), .C(n30332), .Z(n28377)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i21318_2_lut_rep_474 (.A(count[11]), .B(count[10]), .Z(n30483)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21318_2_lut_rep_474.init = 16'heeee;
    LUT4 i21434_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n28587)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21434_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_475 (.A(count[2]), .B(count[1]), .Z(n30484)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_475.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[0]), 
         .D(n30425), .Z(n28146)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.A(count[2]), .B(count[1]), .C(n30485), 
         .D(n30425), .Z(n28226)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut_adj_34.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_35 (.A(count[2]), .B(count[1]), .C(count[4]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_35.init = 16'hf8f8;
    LUT4 i146_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[3]), .Z(n162)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i146_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_476 (.A(count[8]), .B(count[0]), .Z(n30485)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_476.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_36 (.A(count[8]), .B(count[0]), .C(count[1]), 
         .D(count[2]), .Z(n4_adj_47)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut_adj_36.init = 16'h8000;
    LUT4 i21805_4_lut (.A(n54), .B(n28337), .C(n30369), .D(n10), .Z(n28857)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21805_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n30303), .B(n13181), .C(n11), .D(n28587), .Z(n16272)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i4_4_lut (.A(n28226), .B(n28337), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i1_2_lut (.A(count[7]), .B(count[6]), .Z(n20243)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_37 (.A(n1037), .B(n1025), .Z(n28337)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_37.init = 16'hbbbb;
    LUT4 i1_2_lut_adj_38 (.A(count[15]), .B(count[14]), .Z(n13181)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_38.init = 16'heeee;
    LUT4 i2_4_lut_adj_39 (.A(n20243), .B(count[5]), .C(count[3]), .D(n4), 
         .Z(n26341)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_39.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n13181), .D(n30483), 
         .Z(n13179)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(n30425), .B(n28431), .C(n30392), .D(n4_adj_47), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i21284_3_lut (.A(n13179), .B(count[9]), .C(n154), .Z(n28431)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i21284_3_lut.init = 16'heaea;
    LUT4 i15109_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15109_2_lut_4_lut.init = 16'h0400;
    LUT4 i15108_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15108_2_lut_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    CCU2D sub_65_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25826), 
          .S0(n941[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_9.INIT1 = 16'h0000;
    defparam sub_65_add_2_9.INJECT1_0 = "NO";
    defparam sub_65_add_2_9.INJECT1_1 = "NO";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    CCU2D sub_65_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25825), 
          .COUT(n25826), .S0(n941[5]), .S1(n941[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_65_add_2_7.INJECT1_0 = "NO";
    defparam sub_65_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_65_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25824), 
          .COUT(n25825), .S0(n941[3]), .S1(n941[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_65_add_2_5.INJECT1_0 = "NO";
    defparam sub_65_add_2_5.INJECT1_1 = "NO";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D sub_65_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25823), 
          .COUT(n25824), .S0(n941[1]), .S1(n941[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_65_add_2_3.INJECT1_0 = "NO";
    defparam sub_65_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_65_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25823), 
          .S1(n941[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_1.INIT0 = 16'hF000;
    defparam sub_65_add_2_1.INIT1 = 16'h5555;
    defparam sub_65_add_2_1.INJECT1_0 = "NO";
    defparam sub_65_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1752_17 (.A0(count[15]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25562), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_17.INIT0 = 16'hd222;
    defparam add_1752_17.INIT1 = 16'h0000;
    defparam add_1752_17.INJECT1_0 = "NO";
    defparam add_1752_17.INJECT1_1 = "NO";
    CCU2D add_1752_15 (.A0(count[13]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n30482), .C1(GND_net), .D1(GND_net), .CIN(n25561), 
          .COUT(n25562), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_15.INIT0 = 16'hd222;
    defparam add_1752_15.INIT1 = 16'hd222;
    defparam add_1752_15.INJECT1_0 = "NO";
    defparam add_1752_15.INJECT1_1 = "NO";
    CCU2D add_1752_13 (.A0(count[11]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n30482), .C1(GND_net), .D1(GND_net), .CIN(n25560), 
          .COUT(n25561), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_13.INIT0 = 16'hd222;
    defparam add_1752_13.INIT1 = 16'hd222;
    defparam add_1752_13.INJECT1_0 = "NO";
    defparam add_1752_13.INJECT1_1 = "NO";
    LUT4 i15107_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15107_2_lut_4_lut.init = 16'h0400;
    CCU2D add_1752_11 (.A0(count[9]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n30482), .C1(GND_net), .D1(GND_net), .CIN(n25559), 
          .COUT(n25560), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_11.INIT0 = 16'hd222;
    defparam add_1752_11.INIT1 = 16'hd222;
    defparam add_1752_11.INJECT1_0 = "NO";
    defparam add_1752_11.INJECT1_1 = "NO";
    CCU2D add_1752_9 (.A0(count[7]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n30482), .C1(GND_net), .D1(GND_net), .CIN(n25558), 
          .COUT(n25559), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_9.INIT0 = 16'hd222;
    defparam add_1752_9.INIT1 = 16'hd222;
    defparam add_1752_9.INJECT1_0 = "NO";
    defparam add_1752_9.INJECT1_1 = "NO";
    LUT4 i21671_4_lut (.A(n28021), .B(n30482), .C(n30332), .D(n28337), 
         .Z(n28723)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i21671_4_lut.init = 16'h3031;
    LUT4 i2_4_lut_adj_40 (.A(n28020), .B(n30368), .C(n28146), .D(n26341), 
         .Z(n28021)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i2_4_lut_adj_40.init = 16'ha888;
    LUT4 i3_3_lut (.A(n54), .B(n28431), .C(n30369), .Z(n28020)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i3_3_lut.init = 16'h1010;
    LUT4 i2_4_lut_adj_41 (.A(n30483), .B(count[9]), .C(n20243), .D(n4_adj_48), 
         .Z(n28286)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_41.init = 16'hfeee;
    LUT4 i1_4_lut (.A(count[8]), .B(count[4]), .C(n162), .D(count[5]), 
         .Z(n4_adj_48)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut.init = 16'haaa8;
    LUT4 i21780_3_lut_3_lut_4_lut (.A(n26341), .B(n30368), .C(n28431), 
         .D(n30332), .Z(n28378)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i21780_3_lut_3_lut_4_lut.init = 16'h000e;
    CCU2D add_1752_7 (.A0(count[5]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n30482), .C1(GND_net), .D1(GND_net), .CIN(n25557), 
          .COUT(n25558), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_7.INIT0 = 16'hd222;
    defparam add_1752_7.INIT1 = 16'hd222;
    defparam add_1752_7.INJECT1_0 = "NO";
    defparam add_1752_7.INJECT1_1 = "NO";
    LUT4 i15106_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15106_2_lut_4_lut.init = 16'h0400;
    LUT4 i23_4_lut (.A(n30458), .B(count[2]), .C(n30459), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i15105_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15105_2_lut_4_lut.init = 16'h0400;
    LUT4 i15104_2_lut_4_lut (.A(n30392), .B(count[8]), .C(n30393), .D(n941[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15104_2_lut_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14306), .PD(n16272), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX valid_48 (.D(n28378), .SP(n26592), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1031));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D add_1752_5 (.A0(count[3]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n30482), .C1(GND_net), .D1(GND_net), .CIN(n25556), 
          .COUT(n25557), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_5.INIT0 = 16'hd222;
    defparam add_1752_5.INIT1 = 16'hd222;
    defparam add_1752_5.INJECT1_0 = "NO";
    defparam add_1752_5.INJECT1_1 = "NO";
    CCU2D add_1752_3 (.A0(count[1]), .B0(n30482), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n30482), .C1(GND_net), .D1(GND_net), .CIN(n25555), 
          .COUT(n25556), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_3.INIT0 = 16'hd222;
    defparam add_1752_3.INIT1 = 16'hd222;
    defparam add_1752_3.INJECT1_0 = "NO";
    defparam add_1752_3.INJECT1_1 = "NO";
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n30392), .C(n28146), 
         .D(n26341), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    CCU2D add_1752_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28377), .B1(n1037), .C1(count[0]), .D1(n1025), .COUT(n25555), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1752_1.INIT0 = 16'hF000;
    defparam add_1752_1.INIT1 = 16'ha565;
    defparam add_1752_1.INJECT1_0 = "NO";
    defparam add_1752_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (n28855, n30303, debug_c_c, rc_ch3_c, GND_net, 
            n1016, n26607, \register[3] , n14307, n28770) /* synthesis syn_module_defined=1 */ ;
    output n28855;
    input n30303;
    input debug_c_c;
    input rc_ch3_c;
    input GND_net;
    output n1016;
    input n26607;
    output [7:0]\register[3] ;
    input n14307;
    output n28770;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30450, n26703, n30329, n21658, n28307;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n13158, n30381, n30382, n30354, n30355, n26331, n54, 
        n28346, n10, n11, n28583, n16274, n28264, n154, n1022, 
        n1010, n30446, n28308, n152, n103, n30447, n30407, n30448, 
        n6, n4, n4_adj_43, n30449, n30456, n30457, n5, n25570;
    wire [15:0]n116;
    
    wire n25569, n25568;
    wire [7:0]n43;
    
    wire n25830;
    wire [7:0]n932;
    
    wire n25829, n25828, n25827, n25567, n25566, n25565, n25564, 
        n25563, n5_adj_44, n28537, n6_adj_45, n26606, n4_adj_46;
    
    LUT4 i21775_3_lut_3_lut_4_lut (.A(n30450), .B(n26703), .C(n30329), 
         .D(n21658), .Z(n28307)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21775_3_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_372 (.A(count[9]), .B(n13158), .Z(n30381)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_372.init = 16'heeee;
    LUT4 i1_3_lut_rep_345_4_lut (.A(count[9]), .B(n13158), .C(n30382), 
         .D(count[8]), .Z(n30354)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_3_lut_rep_345_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_346_3_lut (.A(count[9]), .B(n13158), .C(count[8]), 
         .Z(n30355)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_346_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_320_3_lut_4_lut (.A(count[9]), .B(n13158), .C(n26331), 
         .D(count[8]), .Z(n30329)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_320_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21803_4_lut (.A(n54), .B(n28346), .C(n30354), .D(n10), .Z(n28855)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21803_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n30303), .B(n30450), .C(n11), .D(n28583), .Z(n16274)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i4_4_lut (.A(n28264), .B(n28346), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n30303), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1022));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i5_2_lut_rep_437 (.A(n1010), .B(n1022), .Z(n30446)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_437.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1010), .B(n1022), .C(n26703), .D(n30450), 
         .Z(n28308)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    PFUMX i13937 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    LUT4 i1_2_lut_rep_438 (.A(count[7]), .B(count[6]), .Z(n30447)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_438.init = 16'h8888;
    LUT4 i1_2_lut_rep_398_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n30407)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_398_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n30448), 
         .D(count[8]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_439 (.A(count[2]), .B(count[1]), .Z(n30448)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_439.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4_adj_43)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i21310_2_lut_rep_440 (.A(count[11]), .B(count[10]), .Z(n30449)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21310_2_lut_rep_440.init = 16'heeee;
    LUT4 i21430_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n28583)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21430_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_441 (.A(count[15]), .B(count[14]), .Z(n30450)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_441.init = 16'heeee;
    LUT4 i2_3_lut_rep_447 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n30456)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_447.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[8]), .D(n30457), 
         .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_448 (.A(count[4]), .B(count[5]), .Z(n30457)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_448.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_28 (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n5)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut_adj_28.init = 16'h8000;
    FD1P3IX valid_48 (.D(n28307), .SP(n26607), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1016));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i3_3_lut_rep_373_4_lut (.A(count[3]), .B(n30457), .C(n30447), 
         .D(n30448), .Z(n30382)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_3_lut_rep_373_4_lut.init = 16'h8000;
    CCU2D add_1748_17 (.A0(count[15]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25570), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_17.INIT0 = 16'hd222;
    defparam add_1748_17.INIT1 = 16'h0000;
    defparam add_1748_17.INJECT1_0 = "NO";
    defparam add_1748_17.INJECT1_1 = "NO";
    FD1P3AX prev_in_46 (.D(n1022), .SP(n30303), .CK(debug_c_c), .Q(n1010));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D add_1748_15 (.A0(count[13]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n30446), .C1(GND_net), .D1(GND_net), .CIN(n25569), 
          .COUT(n25570), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_15.INIT0 = 16'hd222;
    defparam add_1748_15.INIT1 = 16'hd222;
    defparam add_1748_15.INJECT1_0 = "NO";
    defparam add_1748_15.INJECT1_1 = "NO";
    CCU2D add_1748_13 (.A0(count[11]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n30446), .C1(GND_net), .D1(GND_net), .CIN(n25568), 
          .COUT(n25569), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_13.INIT0 = 16'hd222;
    defparam add_1748_13.INIT1 = 16'hd222;
    defparam add_1748_13.INJECT1_0 = "NO";
    defparam add_1748_13.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D sub_64_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25830), 
          .S0(n932[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_9.INIT1 = 16'h0000;
    defparam sub_64_add_2_9.INJECT1_0 = "NO";
    defparam sub_64_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25829), 
          .COUT(n25830), .S0(n932[5]), .S1(n932[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_64_add_2_7.INJECT1_0 = "NO";
    defparam sub_64_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25828), 
          .COUT(n25829), .S0(n932[3]), .S1(n932[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_64_add_2_5.INJECT1_0 = "NO";
    defparam sub_64_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25827), 
          .COUT(n25828), .S0(n932[1]), .S1(n932[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_64_add_2_3.INJECT1_0 = "NO";
    defparam sub_64_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25827), 
          .S1(n932[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_1.INIT0 = 16'hF000;
    defparam sub_64_add_2_1.INIT1 = 16'h5555;
    defparam sub_64_add_2_1.INJECT1_0 = "NO";
    defparam sub_64_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1748_11 (.A0(count[9]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n30446), .C1(GND_net), .D1(GND_net), .CIN(n25567), 
          .COUT(n25568), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_11.INIT0 = 16'hd222;
    defparam add_1748_11.INIT1 = 16'hd222;
    defparam add_1748_11.INJECT1_0 = "NO";
    defparam add_1748_11.INJECT1_1 = "NO";
    CCU2D add_1748_9 (.A0(count[7]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n30446), .C1(GND_net), .D1(GND_net), .CIN(n25566), 
          .COUT(n25567), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_9.INIT0 = 16'hd222;
    defparam add_1748_9.INIT1 = 16'hd222;
    defparam add_1748_9.INJECT1_0 = "NO";
    defparam add_1748_9.INJECT1_1 = "NO";
    CCU2D add_1748_7 (.A0(count[5]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n30446), .C1(GND_net), .D1(GND_net), .CIN(n25565), 
          .COUT(n25566), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_7.INIT0 = 16'hd222;
    defparam add_1748_7.INIT1 = 16'hd222;
    defparam add_1748_7.INJECT1_0 = "NO";
    defparam add_1748_7.INJECT1_1 = "NO";
    CCU2D add_1748_5 (.A0(count[3]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n30446), .C1(GND_net), .D1(GND_net), .CIN(n25564), 
          .COUT(n25565), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_5.INIT0 = 16'hd222;
    defparam add_1748_5.INIT1 = 16'hd222;
    defparam add_1748_5.INJECT1_0 = "NO";
    defparam add_1748_5.INJECT1_1 = "NO";
    CCU2D add_1748_3 (.A0(count[1]), .B0(n30446), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n30446), .C1(GND_net), .D1(GND_net), .CIN(n25563), 
          .COUT(n25564), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_3.INIT0 = 16'hd222;
    defparam add_1748_3.INIT1 = 16'hd222;
    defparam add_1748_3.INJECT1_0 = "NO";
    defparam add_1748_3.INJECT1_1 = "NO";
    CCU2D add_1748_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28308), .B1(n1022), .C1(count[0]), .D1(n1010), .COUT(n25563), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1748_1.INIT0 = 16'hF000;
    defparam add_1748_1.INIT1 = 16'ha565;
    defparam add_1748_1.INJECT1_0 = "NO";
    defparam add_1748_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_29 (.A(n30381), .B(count[8]), .C(n30382), 
         .D(n54), .Z(n5_adj_44)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_29.init = 16'h00fb;
    LUT4 i15102_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15102_2_lut_4_lut.init = 16'h0400;
    LUT4 i15101_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15101_2_lut_4_lut.init = 16'h0400;
    LUT4 i15100_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15100_2_lut_4_lut.init = 16'h0400;
    LUT4 i15099_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15099_2_lut_4_lut.init = 16'h0400;
    LUT4 i15098_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15098_2_lut_4_lut.init = 16'h0400;
    LUT4 i15097_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15097_2_lut_4_lut.init = 16'h0400;
    LUT4 i15096_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15096_2_lut_4_lut.init = 16'h0400;
    LUT4 i14862_2_lut_4_lut (.A(n30381), .B(count[8]), .C(n30382), .D(n932[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14862_2_lut_4_lut.init = 16'h0400;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[0]), .B(n30382), .C(n30355), 
         .D(n26331), .Z(n10)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0700;
    LUT4 i21387_3_lut_4_lut (.A(count[0]), .B(n30382), .C(n26331), .D(n30355), 
         .Z(n28537)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21387_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_3_lut_adj_30 (.A(count[0]), .B(n30382), .C(count[8]), 
         .Z(n28264)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_30.init = 16'h8080;
    LUT4 i23_4_lut (.A(n30456), .B(count[2]), .C(n30457), .D(n6_adj_45), 
         .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6_adj_45)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14307), .PD(n16274), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i21718_4_lut (.A(n30450), .B(n30446), .C(n26703), .D(n26606), 
         .Z(n28770)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i21718_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5_adj_44), .B(n28346), .C(n28537), .D(n21658), 
         .Z(n26606)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i15275_3_lut (.A(count[9]), .B(n13158), .C(n154), .Z(n21658)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15275_3_lut.init = 16'hecec;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n30450), .D(n30449), 
         .Z(n13158)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_31 (.A(n30447), .B(count[5]), .C(count[3]), .D(n4_adj_43), 
         .Z(n26331)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_31.init = 16'h8880;
    LUT4 i2_4_lut_adj_32 (.A(count[13]), .B(count[12]), .C(n30449), .D(n4_adj_46), 
         .Z(n26703)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_32.init = 16'h8880;
    LUT4 i1_4_lut_adj_33 (.A(count[9]), .B(count[4]), .C(n30407), .D(n4), 
         .Z(n4_adj_46)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_33.init = 16'hfaea;
    LUT4 i21_4_lut (.A(n5), .B(n21658), .C(n30381), .D(n6), .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_2_lut (.A(n1022), .B(n1010), .Z(n28346)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (GND_net, n28853, n30303, n1001, debug_c_c, 
            n26604, \register[2] , n14308, rc_ch2_c, n28773) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n28853;
    input n30303;
    output n1001;
    input debug_c_c;
    input n26604;
    output [7:0]\register[2] ;
    input n14308;
    input rc_ch2_c;
    output n28773;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25575;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n5;
    wire [15:0]n116;
    
    wire n25576, n25574, n30336, n28439, n30335, n26322, n28313, 
        n54, n28340, n30333, n10, n30412, n16, n16276, n26, 
        n30386, n154, n30466, n30360, n5_adj_40;
    wire [7:0]n923;
    wire [7:0]n43;
    
    wire n25573, n25572, n28355, n28140, n28539, n152, n103, n25571, 
        n995, n1007, n30455, n30468, n28314, n30467, n26772, n20429, 
        n30414, n30469, n4, n4_adj_41, n30384, n25834, n25833, 
        n25832, n25831, n26603, n4_adj_42, n26501, n6, n25578, 
        n25577;
    
    CCU2D add_1744_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25575), 
          .COUT(n25576), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_11.INIT0 = 16'hd222;
    defparam add_1744_11.INIT1 = 16'hd222;
    defparam add_1744_11.INJECT1_0 = "NO";
    defparam add_1744_11.INJECT1_1 = "NO";
    CCU2D add_1744_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25574), 
          .COUT(n25575), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_9.INIT0 = 16'hd222;
    defparam add_1744_9.INIT1 = 16'hd222;
    defparam add_1744_9.INJECT1_0 = "NO";
    defparam add_1744_9.INJECT1_1 = "NO";
    LUT4 i21771_3_lut_4_lut_4_lut (.A(n30336), .B(n28439), .C(n30335), 
         .D(n26322), .Z(n28313)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i21771_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i21801_4_lut (.A(n54), .B(n28340), .C(n30333), .D(n10), .Z(n28853)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21801_4_lut.init = 16'h3323;
    LUT4 i8_4_lut (.A(n30412), .B(n16), .C(count[13]), .D(count[11]), 
         .Z(n16276)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i8_4_lut.init = 16'h0004;
    LUT4 i7_4_lut (.A(count[10]), .B(n30303), .C(n26), .D(n28340), .Z(n16)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i7_4_lut.init = 16'h0040;
    LUT4 i33_4_lut (.A(n30386), .B(n154), .C(count[9]), .D(n30466), 
         .Z(n26)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_4_lut.init = 16'h3a30;
    LUT4 i1_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n54), 
         .Z(n5_adj_40)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h00fb;
    LUT4 i15090_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15090_2_lut_4_lut.init = 16'h0400;
    LUT4 i15089_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15089_2_lut_4_lut.init = 16'h0400;
    LUT4 i15088_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15088_2_lut_4_lut.init = 16'h0400;
    FD1P3IX valid_48 (.D(n28313), .SP(n26604), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1001));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D add_1744_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25573), 
          .COUT(n25574), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_7.INIT0 = 16'hd222;
    defparam add_1744_7.INIT1 = 16'hd222;
    defparam add_1744_7.INJECT1_0 = "NO";
    defparam add_1744_7.INJECT1_1 = "NO";
    CCU2D add_1744_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25572), 
          .COUT(n25573), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_5.INIT0 = 16'hd222;
    defparam add_1744_5.INIT1 = 16'hd222;
    defparam add_1744_5.INJECT1_0 = "NO";
    defparam add_1744_5.INJECT1_1 = "NO";
    LUT4 i15087_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15087_2_lut_4_lut.init = 16'h0400;
    LUT4 i15086_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15086_2_lut_4_lut.init = 16'h0400;
    LUT4 i15085_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15085_2_lut_4_lut.init = 16'h0400;
    LUT4 i15084_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15084_2_lut_4_lut.init = 16'h0400;
    LUT4 i14855_2_lut_4_lut (.A(n30360), .B(count[8]), .C(n30386), .D(n923[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14855_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_351_4_lut (.A(n30412), .B(count[13]), .C(n28355), 
         .D(count[9]), .Z(n30360)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_351_4_lut.init = 16'hfffe;
    LUT4 i21388_3_lut_4_lut (.A(count[8]), .B(n30360), .C(n26322), .D(n28140), 
         .Z(n28539)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i21388_3_lut_4_lut.init = 16'hfeee;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n30360), .C(n28140), 
         .D(n26322), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    PFUMX i14031 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    CCU2D add_1744_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25571), 
          .COUT(n25572), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_3.INIT0 = 16'hd222;
    defparam add_1744_3.INIT1 = 16'hd222;
    defparam add_1744_3.INJECT1_0 = "NO";
    defparam add_1744_3.INJECT1_1 = "NO";
    LUT4 i5_2_lut (.A(n995), .B(n1007), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_rep_446 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n30455)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_446.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_20 (.A(count[7]), .B(count[6]), .C(count[8]), 
         .D(n30468), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_20.init = 16'hfffe;
    CCU2D add_1744_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28314), .B1(n1007), .C1(count[0]), .D1(n995), .COUT(n25571), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_1.INIT0 = 16'hF000;
    defparam add_1744_1.INIT1 = 16'ha565;
    defparam add_1744_1.INJECT1_0 = "NO";
    defparam add_1744_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_457 (.A(count[8]), .B(count[0]), .Z(n30466)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_457.init = 16'h8888;
    LUT4 i1_2_lut_rep_458 (.A(count[15]), .B(count[14]), .Z(n30467)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_458.init = 16'heeee;
    LUT4 i1_2_lut_rep_327_3_lut (.A(count[15]), .B(count[14]), .C(n26772), 
         .Z(n30336)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_327_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n26772), 
         .Z(n28314)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21290_2_lut_rep_403_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n30412)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i21290_2_lut_rep_403_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_459 (.A(count[4]), .B(count[5]), .Z(n30468)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_459.init = 16'h8888;
    LUT4 i1_3_lut_rep_405_4_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .D(n20429), .Z(n30414)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_rep_405_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_460 (.A(count[2]), .B(count[1]), .Z(n30469)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_460.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_21 (.A(count[2]), .B(count[1]), .C(count[0]), 
         .D(n30414), .Z(n28140)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut_adj_21.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_22 (.A(count[2]), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n4_adj_41)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut_adj_22.init = 16'h8000;
    LUT4 i3_3_lut_rep_375_4_lut (.A(count[12]), .B(n30467), .C(n28355), 
         .D(count[13]), .Z(n30384)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_375_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_rep_377_4_lut (.A(n20429), .B(count[3]), .C(n30468), 
         .D(n30469), .Z(n30386)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut_rep_377_4_lut.init = 16'h8000;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    CCU2D sub_63_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25834), 
          .S0(n923[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_9.INIT1 = 16'h0000;
    defparam sub_63_add_2_9.INJECT1_0 = "NO";
    defparam sub_63_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25833), 
          .COUT(n25834), .S0(n923[5]), .S1(n923[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_63_add_2_7.INJECT1_0 = "NO";
    defparam sub_63_add_2_7.INJECT1_1 = "NO";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D sub_63_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25832), 
          .COUT(n25833), .S0(n923[3]), .S1(n923[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_63_add_2_5.INJECT1_0 = "NO";
    defparam sub_63_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25831), 
          .COUT(n25832), .S0(n923[1]), .S1(n923[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_63_add_2_3.INJECT1_0 = "NO";
    defparam sub_63_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25831), 
          .S1(n923[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_1.INIT0 = 16'hF000;
    defparam sub_63_add_2_1.INIT1 = 16'h5555;
    defparam sub_63_add_2_1.INJECT1_0 = "NO";
    defparam sub_63_add_2_1.INJECT1_1 = "NO";
    FD1P3AX prev_in_46 (.D(n1007), .SP(n30303), .CK(debug_c_c), .Q(n995));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n30303), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1007));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i21721_4_lut (.A(n30467), .B(n5), .C(n26772), .D(n26603), .Z(n28773)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i21721_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5_adj_40), .B(n28340), .C(n28539), .D(n28439), 
         .Z(n26603)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i2_4_lut (.A(n20429), .B(count[5]), .C(count[3]), .D(n4), .Z(n26322)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_2_lut (.A(count[7]), .B(count[6]), .Z(n20429)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_23 (.A(count[10]), .B(count[11]), .Z(n28355)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_23.init = 16'heeee;
    LUT4 i21_4_lut (.A(n30414), .B(n28439), .C(n30360), .D(n4_adj_41), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i21292_3_lut (.A(n30384), .B(count[9]), .C(n154), .Z(n28439)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i21292_3_lut.init = 16'heaea;
    LUT4 i1_2_lut_adj_24 (.A(n1007), .B(n995), .Z(n28340)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_24.init = 16'hbbbb;
    LUT4 i2_4_lut_adj_25 (.A(count[13]), .B(count[12]), .C(n28355), .D(n4_adj_42), 
         .Z(n26772)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_25.init = 16'h8880;
    LUT4 i1_4_lut_adj_26 (.A(count[9]), .B(n20429), .C(count[8]), .D(n26501), 
         .Z(n4_adj_42)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_26.init = 16'heaaa;
    LUT4 i2_4_lut_adj_27 (.A(count[4]), .B(count[3]), .C(count[5]), .D(n30469), 
         .Z(n26501)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_27.init = 16'hfefa;
    LUT4 i2_3_lut_rep_324_4_lut (.A(count[9]), .B(n30384), .C(n30386), 
         .D(count[8]), .Z(n30333)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i2_3_lut_rep_324_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_326_3_lut (.A(count[9]), .B(n30384), .C(count[8]), 
         .Z(n30335)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_326_3_lut.init = 16'hfefe;
    LUT4 i23_4_lut (.A(n30455), .B(count[2]), .C(n30468), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14308), .PD(n16276), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1744_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25578), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_17.INIT0 = 16'hd222;
    defparam add_1744_17.INIT1 = 16'h0000;
    defparam add_1744_17.INJECT1_0 = "NO";
    defparam add_1744_17.INJECT1_1 = "NO";
    CCU2D add_1744_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25577), 
          .COUT(n25578), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_15.INIT0 = 16'hd222;
    defparam add_1744_15.INIT1 = 16'hd222;
    defparam add_1744_15.INJECT1_0 = "NO";
    defparam add_1744_15.INJECT1_1 = "NO";
    CCU2D add_1744_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n25576), 
          .COUT(n25577), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1744_13.INIT0 = 16'hd222;
    defparam add_1744_13.INIT1 = 16'hd222;
    defparam add_1744_13.INJECT1_0 = "NO";
    defparam add_1744_13.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (debug_c_c, n30303, GND_net, n32380, n28851, 
            \register[1] , n14309, rc_ch1_c, n28725, n986, n26596) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n30303;
    input GND_net;
    input n32380;
    output n28851;
    output [7:0]\register[1] ;
    input n14309;
    input rc_ch1_c;
    output n28725;
    output n986;
    input n26596;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n30428, n30399, n30429, n28252, n28182, n30347, n28486, 
        n30334, n28372, n4, n13118, n5, n6, n26493, n13207, 
        n28297;
    wire [7:0]n914;
    
    wire n23;
    wire [7:0]n43;
    wire [15:0]n116;
    
    wire n980, n992, n28299, n30397, n30348, n21674, n30346, n30474, 
        n28371, n115, n30490, n26656, n18, n28042, n30320, n28496, 
        n30319, n25838, n25837, n16278, n25836, n25835, n25586, 
        n25585, n25584, n25583, n28241, n4_adj_39, n25582, n25581, 
        n25580, n25579;
    
    LUT4 i1_2_lut_rep_419 (.A(count[7]), .B(count[6]), .Z(n30428)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_419.init = 16'h8888;
    LUT4 i1_2_lut_rep_390_3_lut (.A(count[7]), .B(count[6]), .C(count[5]), 
         .Z(n30399)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_390_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_420 (.A(count[2]), .B(count[3]), .Z(n30429)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_420.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n28252)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i21769_3_lut_3_lut_4_lut (.A(n28182), .B(n30347), .C(n28486), 
         .D(n30334), .Z(n28372)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i21769_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_4_lut (.A(count[2]), .B(n30399), .C(n4), .D(count[1]), .Z(n28182)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut.init = 16'hc8c0;
    LUT4 i1_2_lut (.A(count[4]), .B(count[3]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i21339_4_lut (.A(n13118), .B(count[9]), .C(n5), .D(n6), .Z(n28486)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i21339_4_lut.init = 16'heeea;
    LUT4 i1_4_lut_adj_9 (.A(count[6]), .B(count[5]), .C(n26493), .D(count[4]), 
         .Z(n5)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_9.init = 16'heaaa;
    LUT4 i2_2_lut (.A(count[7]), .B(count[8]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(count[2]), .B(count[1]), .C(count[0]), .D(count[3]), 
         .Z(n26493)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_10 (.A(count[12]), .B(count[13]), .C(n13207), .D(n28297), 
         .Z(n13118)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_10.init = 16'hfffe;
    LUT4 i1_2_lut_adj_11 (.A(count[15]), .B(count[14]), .Z(n13207)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_11.init = 16'heeee;
    LUT4 i1_2_lut_adj_12 (.A(count[11]), .B(count[10]), .Z(n28297)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_12.init = 16'heeee;
    LUT4 i15074_2_lut (.A(n914[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15074_2_lut.init = 16'h8888;
    LUT4 i15073_2_lut (.A(n914[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15073_2_lut.init = 16'h8888;
    LUT4 i15072_2_lut (.A(n914[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15072_2_lut.init = 16'h8888;
    LUT4 i15071_2_lut (.A(n914[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15071_2_lut.init = 16'h8888;
    LUT4 i15070_2_lut (.A(n914[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15070_2_lut.init = 16'h8888;
    LUT4 i15069_2_lut (.A(n914[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15069_2_lut.init = 16'h8888;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n992), .SP(n30303), .CK(debug_c_c), .Q(n980));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_4_lut_rep_325 (.A(n13207), .B(count[13]), .C(count[12]), .D(n28299), 
         .Z(n30334)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_325.init = 16'heaaa;
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_388 (.A(count[9]), .B(n13118), .Z(n30397)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_388.init = 16'heeee;
    LUT4 i1_2_lut_rep_338_3_lut (.A(count[9]), .B(n13118), .C(count[8]), 
         .Z(n30347)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_338_3_lut.init = 16'hfefe;
    LUT4 i15290_2_lut_3_lut_4_lut (.A(count[9]), .B(n13118), .C(n30348), 
         .D(count[8]), .Z(n21674)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i15290_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_337_3_lut_4_lut (.A(count[9]), .B(n13118), .C(n28182), 
         .D(count[8]), .Z(n30346)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_337_3_lut_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut_rep_465 (.A(n980), .B(n992), .Z(n30474)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_465.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_13 (.A(n980), .B(n992), .C(n30334), .Z(n28371)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_adj_13.init = 16'hf4f4;
    LUT4 i2_3_lut_4_lut (.A(count[5]), .B(n30428), .C(count[4]), .D(n30429), 
         .Z(n115)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_481 (.A(n992), .B(n980), .Z(n30490)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_481.init = 16'hbbbb;
    LUT4 i3_4_lut_adj_14 (.A(n26656), .B(n992), .C(n32380), .D(n18), 
         .Z(n28042)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_14.init = 16'h0200;
    LUT4 i21799_2_lut_3_lut (.A(n992), .B(n980), .C(n26656), .Z(n28851)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i21799_2_lut_3_lut.init = 16'h4040;
    LUT4 i21349_3_lut_4_lut (.A(n30320), .B(n28486), .C(n30397), .D(n23), 
         .Z(n28496)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21349_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21_3_lut_rep_310_4_lut (.A(count[8]), .B(n30348), .C(n30397), 
         .D(n28486), .Z(n30319)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21_3_lut_rep_310_4_lut.init = 16'h00f8;
    LUT4 i1_2_lut_3_lut_adj_15 (.A(count[8]), .B(n30348), .C(count[9]), 
         .Z(n18)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_15.init = 16'hf8f8;
    CCU2D sub_62_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25838), 
          .S0(n914[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_9.INIT1 = 16'h0000;
    defparam sub_62_add_2_9.INJECT1_0 = "NO";
    defparam sub_62_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_62_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25837), 
          .COUT(n25838), .S0(n914[5]), .S1(n914[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_62_add_2_7.INJECT1_0 = "NO";
    defparam sub_62_add_2_7.INJECT1_1 = "NO";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D sub_62_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25836), 
          .COUT(n25837), .S0(n914[3]), .S1(n914[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_62_add_2_5.INJECT1_0 = "NO";
    defparam sub_62_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_62_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25835), 
          .COUT(n25836), .S0(n914[1]), .S1(n914[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_62_add_2_3.INJECT1_0 = "NO";
    defparam sub_62_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_62_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25835), 
          .S1(n914[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_1.INIT0 = 16'hF000;
    defparam sub_62_add_2_1.INIT1 = 16'h5555;
    defparam sub_62_add_2_1.INJECT1_0 = "NO";
    defparam sub_62_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_339 (.A(n115), .B(count[1]), .C(count[0]), .Z(n30348)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_3_lut_rep_339.init = 16'h8080;
    LUT4 i1_2_lut_rep_311_4_lut (.A(n115), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n30320)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_311_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n30303), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n992));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    CCU2D add_1740_17 (.A0(count[15]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25586), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_17.INIT0 = 16'hd222;
    defparam add_1740_17.INIT1 = 16'h0000;
    defparam add_1740_17.INJECT1_0 = "NO";
    defparam add_1740_17.INJECT1_1 = "NO";
    CCU2D add_1740_15 (.A0(count[13]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n30474), .C1(GND_net), .D1(GND_net), .CIN(n25585), 
          .COUT(n25586), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_15.INIT0 = 16'hd222;
    defparam add_1740_15.INIT1 = 16'hd222;
    defparam add_1740_15.INJECT1_0 = "NO";
    defparam add_1740_15.INJECT1_1 = "NO";
    LUT4 i14850_2_lut (.A(n914[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i14850_2_lut.init = 16'h8888;
    CCU2D add_1740_13 (.A0(count[11]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n30474), .C1(GND_net), .D1(GND_net), .CIN(n25584), 
          .COUT(n25585), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_13.INIT0 = 16'hd222;
    defparam add_1740_13.INIT1 = 16'hd222;
    defparam add_1740_13.INJECT1_0 = "NO";
    defparam add_1740_13.INJECT1_1 = "NO";
    CCU2D add_1740_11 (.A0(count[9]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n30474), .C1(GND_net), .D1(GND_net), .CIN(n25583), 
          .COUT(n25584), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_11.INIT0 = 16'hd222;
    defparam add_1740_11.INIT1 = 16'hd222;
    defparam add_1740_11.INJECT1_0 = "NO";
    defparam add_1740_11.INJECT1_1 = "NO";
    LUT4 i21673_4_lut (.A(n28241), .B(n30474), .C(n30334), .D(n30490), 
         .Z(n28725)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i21673_4_lut.init = 16'h3031;
    LUT4 i4_4_lut (.A(n30347), .B(n28496), .C(n30348), .D(n28182), .Z(n28241)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i4_4_lut.init = 16'h3222;
    LUT4 i2_4_lut (.A(n28297), .B(count[9]), .C(count[8]), .D(n4_adj_39), 
         .Z(n28299)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut.init = 16'hfeee;
    LUT4 i1_4_lut_adj_16 (.A(n30428), .B(count[4]), .C(count[5]), .D(n28252), 
         .Z(n4_adj_39)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_16.init = 16'haaa8;
    CCU2D add_1740_9 (.A0(count[7]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n30474), .C1(GND_net), .D1(GND_net), .CIN(n25582), 
          .COUT(n25583), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_9.INIT0 = 16'hd222;
    defparam add_1740_9.INIT1 = 16'hd222;
    defparam add_1740_9.INJECT1_0 = "NO";
    defparam add_1740_9.INJECT1_1 = "NO";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    LUT4 i15075_2_lut (.A(n914[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15075_2_lut.init = 16'h8888;
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_17 (.A(count[8]), .B(n30397), .C(count[1]), .D(n115), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_17.init = 16'h0222;
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_18 (.A(n30319), .B(n23), .C(n30346), .D(n21674), 
         .Z(n26656)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_18.init = 16'heefe;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14309), .PD(n16278), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n30303), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n30303), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    CCU2D add_1740_7 (.A0(count[5]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n30474), .C1(GND_net), .D1(GND_net), .CIN(n25581), 
          .COUT(n25582), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_7.INIT0 = 16'hd222;
    defparam add_1740_7.INIT1 = 16'hd222;
    defparam add_1740_7.INJECT1_0 = "NO";
    defparam add_1740_7.INJECT1_1 = "NO";
    FD1P3IX valid_48 (.D(n28372), .SP(n26596), .CD(GND_net), .CK(debug_c_c), 
            .Q(n986));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D add_1740_5 (.A0(count[3]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n30474), .C1(GND_net), .D1(GND_net), .CIN(n25580), 
          .COUT(n25581), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_5.INIT0 = 16'hd222;
    defparam add_1740_5.INIT1 = 16'hd222;
    defparam add_1740_5.INJECT1_0 = "NO";
    defparam add_1740_5.INJECT1_1 = "NO";
    CCU2D add_1740_3 (.A0(count[1]), .B0(n30474), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n30474), .C1(GND_net), .D1(GND_net), .CIN(n25579), 
          .COUT(n25580), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_3.INIT0 = 16'hd222;
    defparam add_1740_3.INIT1 = 16'hd222;
    defparam add_1740_3.INJECT1_0 = "NO";
    defparam add_1740_3.INJECT1_1 = "NO";
    CCU2D add_1740_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28371), .B1(n992), .C1(count[0]), .D1(n980), .COUT(n25579), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_1.INIT0 = 16'hF000;
    defparam add_1740_1.INIT1 = 16'ha565;
    defparam add_1740_1.INJECT1_0 = "NO";
    defparam add_1740_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_19 (.A(n30303), .B(n28042), .C(n980), .D(n28486), 
         .Z(n16278)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_19.init = 16'h0080;
    
endmodule
//
// Verilog Description of module EncoderPeripheral
//

module EncoderPeripheral (read_value, debug_c_c, n13589, n30321, \read_size[2] , 
            n30380, \register_addr[0] , \read_size[0] , n30370, prev_select, 
            n30361, encoder_ra_c, encoder_rb_c, encoder_ri_c, \register_addr[1] , 
            n30489, n30491, n13269, n30422, n30366, n302, n97, 
            n49, n47, n39, n37, n14013, qreset, \quadA_delayed[1] , 
            GND_net, n6, \register[1][0] , VCC_net, \register[1][24] , 
            \register[1][25] , \register[1][29] , \register[1][30] , \quadB_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n13589;
    input n30321;
    output \read_size[2] ;
    input n30380;
    input \register_addr[0] ;
    output \read_size[0] ;
    input n30370;
    output prev_select;
    input n30361;
    input encoder_ra_c;
    input encoder_rb_c;
    input encoder_ri_c;
    input \register_addr[1] ;
    input n30489;
    input n30491;
    output n13269;
    input n30422;
    output n30366;
    output n302;
    input n97;
    input n49;
    input n47;
    input n39;
    input n37;
    input n14013;
    input qreset;
    output \quadA_delayed[1] ;
    input GND_net;
    output n6;
    output \register[1][0] ;
    input VCC_net;
    output \register[1][24] ;
    output \register[1][25] ;
    output \register[1][29] ;
    output \register[1][30] ;
    output \quadB_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]n180;
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    FD1P3IX read_value__i31 (.D(n180[31]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n180[28]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n180[27]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n180[26]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n180[23]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n180[22]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n180[21]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n180[20]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n180[19]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n180[18]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n180[17]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n180[16]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n180[15]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n180[14]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n180[13]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n180[12]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n180[11]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n180[10]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n180[9]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n180[8]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n180[7]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n180[6]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n180[5]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n180[4]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n180[3]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n180[2]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n180[1]), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_size__i2 (.D(n30380), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i14741_2_lut (.A(\register[1] [19]), .B(\register_addr[0] ), .Z(n180[19])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14741_2_lut.init = 16'h8888;
    FD1P3IX read_size__i1 (.D(n30370), .SP(n13589), .CD(n30321), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i14742_2_lut (.A(\register[1] [18]), .B(\register_addr[0] ), .Z(n180[18])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14742_2_lut.init = 16'h8888;
    FD1S3AX prev_select_126 (.D(n30361), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam prev_select_126.GSR = "ENABLED";
    LUT4 i14743_2_lut (.A(\register[1] [17]), .B(\register_addr[0] ), .Z(n180[17])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14743_2_lut.init = 16'h8888;
    LUT4 i14744_2_lut (.A(\register[1] [16]), .B(\register_addr[0] ), .Z(n180[16])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14744_2_lut.init = 16'h8888;
    LUT4 i14745_2_lut (.A(\register[1] [15]), .B(\register_addr[0] ), .Z(n180[15])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14745_2_lut.init = 16'h8888;
    LUT4 i14746_2_lut (.A(\register[1] [14]), .B(\register_addr[0] ), .Z(n180[14])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14746_2_lut.init = 16'h8888;
    LUT4 i14747_2_lut (.A(\register[1] [13]), .B(\register_addr[0] ), .Z(n180[13])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14747_2_lut.init = 16'h8888;
    LUT4 i14748_2_lut (.A(\register[1] [12]), .B(\register_addr[0] ), .Z(n180[12])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14748_2_lut.init = 16'h8888;
    LUT4 i14749_2_lut (.A(\register[1] [11]), .B(\register_addr[0] ), .Z(n180[11])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14749_2_lut.init = 16'h8888;
    LUT4 i14750_2_lut (.A(\register[1] [10]), .B(\register_addr[0] ), .Z(n180[10])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14750_2_lut.init = 16'h8888;
    LUT4 i14751_2_lut (.A(\register[1] [9]), .B(\register_addr[0] ), .Z(n180[9])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14751_2_lut.init = 16'h8888;
    LUT4 i14752_2_lut (.A(\register[1] [8]), .B(\register_addr[0] ), .Z(n180[8])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14752_2_lut.init = 16'h8888;
    LUT4 i14753_2_lut (.A(\register[1] [7]), .B(\register_addr[0] ), .Z(n180[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14753_2_lut.init = 16'h8888;
    LUT4 i14754_2_lut (.A(\register[1] [6]), .B(\register_addr[0] ), .Z(n180[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14754_2_lut.init = 16'h8888;
    LUT4 i14755_2_lut (.A(\register[1] [5]), .B(\register_addr[0] ), .Z(n180[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14755_2_lut.init = 16'h8888;
    LUT4 i14756_2_lut (.A(\register[1] [4]), .B(\register_addr[0] ), .Z(n180[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14756_2_lut.init = 16'h8888;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_ra_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n180[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_rb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n180[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_ri_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n180[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n30489), .C(n30491), 
         .D(\register_addr[0] ), .Z(n13269)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(78[9:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 equal_138_i15_2_lut_rep_357_3_lut_4_lut (.A(\register_addr[1] ), 
         .B(n30489), .C(n30422), .D(\register_addr[0] ), .Z(n30366)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(78[9:33])
    defparam equal_138_i15_2_lut_rep_357_3_lut_4_lut.init = 16'hfffe;
    LUT4 equal_138_i16_1_lut_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n30489), 
         .C(n30422), .D(\register_addr[0] ), .Z(n302)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(78[9:33])
    defparam equal_138_i16_1_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i14739_2_lut (.A(\register[1] [21]), .B(\register_addr[0] ), .Z(n180[21])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14739_2_lut.init = 16'h8888;
    LUT4 i14740_2_lut (.A(\register[1] [20]), .B(\register_addr[0] ), .Z(n180[20])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14740_2_lut.init = 16'h8888;
    FD1P3AX read_value__i0 (.D(n97), .SP(n13589), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n49), .SP(n13589), .CK(debug_c_c), .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n47), .SP(n13589), .CK(debug_c_c), .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n39), .SP(n13589), .CK(debug_c_c), .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n37), .SP(n13589), .CK(debug_c_c), .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=660, LSE_RLINE=670 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i30.GSR = "ENABLED";
    LUT4 i14733_2_lut (.A(\register[1] [31]), .B(\register_addr[0] ), .Z(n180[31])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14733_2_lut.init = 16'h8888;
    LUT4 i14734_2_lut (.A(\register[1] [28]), .B(\register_addr[0] ), .Z(n180[28])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14734_2_lut.init = 16'h8888;
    LUT4 i14735_2_lut (.A(\register[1] [27]), .B(\register_addr[0] ), .Z(n180[27])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14735_2_lut.init = 16'h8888;
    LUT4 i14736_2_lut (.A(\register[1] [26]), .B(\register_addr[0] ), .Z(n180[26])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14736_2_lut.init = 16'h8888;
    LUT4 i14737_2_lut (.A(\register[1] [23]), .B(\register_addr[0] ), .Z(n180[23])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14737_2_lut.init = 16'h8888;
    LUT4 i14738_2_lut (.A(\register[1] [22]), .B(\register_addr[0] ), .Z(n180[22])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14738_2_lut.init = 16'h8888;
    QuadratureDecoder q (.debug_c_c(debug_c_c), .n14013(n14013), .qreset(qreset), 
            .quadA_delayed({Open_9, \quadA_delayed[1] , Open_10}), .GND_net(GND_net), 
            .n6(n6), .\register[1] ({\register[1] [31], \register[1][30] , 
            \register[1][29] , \register[1] [28:26], \register[1][25] , 
            \register[1][24] , \register[1] [23:1], \register[1][0] }), 
            .VCC_net(VCC_net), .encoder_rb_c(encoder_rb_c), .encoder_ra_c(encoder_ra_c), 
            .\quadB_delayed[1] (\quadB_delayed[1] )) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(93[20] 97[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder
//

module QuadratureDecoder (debug_c_c, n14013, qreset, quadA_delayed, 
            GND_net, n6, \register[1] , VCC_net, encoder_rb_c, encoder_ra_c, 
            \quadB_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n14013;
    input qreset;
    output [2:0]quadA_delayed;
    input GND_net;
    output n6;
    output [31:0]\register[1] ;
    input VCC_net;
    input encoder_rb_c;
    input encoder_ra_c;
    output \quadB_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [31:0]n4156;
    
    wire n26216;
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n26217, n26215, n26214, n26213, n26212, n26211, n26210, 
        n26209, n26208, n26207, n26206, n26205, n26204, n26203, 
        n26202;
    wire [2:0]quadA_delayed_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    FD1P3IX count__i13 (.D(n4156[13]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    CCU2D add_1649_31 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n26216), .COUT(n26217), 
          .S0(n4156[28]), .S1(n4156[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_31.INIT0 = 16'h6969;
    defparam add_1649_31.INIT1 = 16'h6969;
    defparam add_1649_31.INJECT1_0 = "NO";
    defparam add_1649_31.INJECT1_1 = "NO";
    CCU2D add_1649_29 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n26215), .COUT(n26216), 
          .S0(n4156[26]), .S1(n4156[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_29.INIT0 = 16'h6969;
    defparam add_1649_29.INIT1 = 16'h6969;
    defparam add_1649_29.INJECT1_0 = "NO";
    defparam add_1649_29.INJECT1_1 = "NO";
    CCU2D add_1649_27 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n26214), .COUT(n26215), 
          .S0(n4156[24]), .S1(n4156[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_27.INIT0 = 16'h6969;
    defparam add_1649_27.INIT1 = 16'h6969;
    defparam add_1649_27.INJECT1_0 = "NO";
    defparam add_1649_27.INJECT1_1 = "NO";
    CCU2D add_1649_25 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n26213), .COUT(n26214), 
          .S0(n4156[22]), .S1(n4156[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_25.INIT0 = 16'h6969;
    defparam add_1649_25.INIT1 = 16'h6969;
    defparam add_1649_25.INJECT1_0 = "NO";
    defparam add_1649_25.INJECT1_1 = "NO";
    CCU2D add_1649_23 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n26212), .COUT(n26213), 
          .S0(n4156[20]), .S1(n4156[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_23.INIT0 = 16'h6969;
    defparam add_1649_23.INIT1 = 16'h6969;
    defparam add_1649_23.INJECT1_0 = "NO";
    defparam add_1649_23.INJECT1_1 = "NO";
    CCU2D add_1649_21 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n26211), .COUT(n26212), 
          .S0(n4156[18]), .S1(n4156[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_21.INIT0 = 16'h6969;
    defparam add_1649_21.INIT1 = 16'h6969;
    defparam add_1649_21.INJECT1_0 = "NO";
    defparam add_1649_21.INJECT1_1 = "NO";
    CCU2D add_1649_19 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n26210), .COUT(n26211), 
          .S0(n4156[16]), .S1(n4156[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_19.INIT0 = 16'h6969;
    defparam add_1649_19.INIT1 = 16'h6969;
    defparam add_1649_19.INJECT1_0 = "NO";
    defparam add_1649_19.INJECT1_1 = "NO";
    FD1P3IX count__i14 (.D(n4156[14]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    CCU2D add_1649_17 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n26209), .COUT(n26210), 
          .S0(n4156[14]), .S1(n4156[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_17.INIT0 = 16'h6969;
    defparam add_1649_17.INIT1 = 16'h6969;
    defparam add_1649_17.INJECT1_0 = "NO";
    defparam add_1649_17.INJECT1_1 = "NO";
    CCU2D add_1649_15 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n26208), .COUT(n26209), 
          .S0(n4156[12]), .S1(n4156[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_15.INIT0 = 16'h6969;
    defparam add_1649_15.INIT1 = 16'h6969;
    defparam add_1649_15.INJECT1_0 = "NO";
    defparam add_1649_15.INJECT1_1 = "NO";
    CCU2D add_1649_13 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n26207), .COUT(n26208), 
          .S0(n4156[10]), .S1(n4156[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_13.INIT0 = 16'h6969;
    defparam add_1649_13.INIT1 = 16'h6969;
    defparam add_1649_13.INJECT1_0 = "NO";
    defparam add_1649_13.INJECT1_1 = "NO";
    CCU2D add_1649_11 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n26206), .COUT(n26207), 
          .S0(n4156[8]), .S1(n4156[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_11.INIT0 = 16'h6969;
    defparam add_1649_11.INIT1 = 16'h6969;
    defparam add_1649_11.INJECT1_0 = "NO";
    defparam add_1649_11.INJECT1_1 = "NO";
    CCU2D add_1649_9 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n26205), .COUT(n26206), 
          .S0(n4156[6]), .S1(n4156[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_9.INIT0 = 16'h6969;
    defparam add_1649_9.INIT1 = 16'h6969;
    defparam add_1649_9.INJECT1_0 = "NO";
    defparam add_1649_9.INJECT1_1 = "NO";
    CCU2D add_1649_7 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n26204), .COUT(n26205), 
          .S0(n4156[4]), .S1(n4156[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_7.INIT0 = 16'h6969;
    defparam add_1649_7.INIT1 = 16'h6969;
    defparam add_1649_7.INJECT1_0 = "NO";
    defparam add_1649_7.INJECT1_1 = "NO";
    FD1P3IX count__i15 (.D(n4156[15]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n4156[16]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n4156[17]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    CCU2D add_1649_5 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n26203), .COUT(n26204), 
          .S0(n4156[2]), .S1(n4156[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_5.INIT0 = 16'h6969;
    defparam add_1649_5.INIT1 = 16'h6969;
    defparam add_1649_5.INJECT1_0 = "NO";
    defparam add_1649_5.INJECT1_1 = "NO";
    CCU2D add_1649_3 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n26202), .COUT(n26203), 
          .S0(n4156[0]), .S1(n4156[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_3.INIT0 = 16'h9696;
    defparam add_1649_3.INIT1 = 16'h6969;
    defparam add_1649_3.INJECT1_0 = "NO";
    defparam add_1649_3.INJECT1_1 = "NO";
    CCU2D add_1649_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26202));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_1.INIT0 = 16'hF000;
    defparam add_1649_1.INIT1 = 16'h6666;
    defparam add_1649_1.INJECT1_0 = "NO";
    defparam add_1649_1.INJECT1_1 = "NO";
    FD1P3IX count__i18 (.D(n4156[18]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n4156[19]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n4156[20]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n4156[21]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n4156[22]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n4156[23]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n4156[24]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n4156[25]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n4156[26]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n4156[27]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n4156[28]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n4156[29]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4156[30]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i31 (.D(n4156[31]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed_c[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_rb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_ra_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed_c[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    FD1P3IX count__i0 (.D(n4156[0]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n4156[1]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n4156[2]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed_c[0]), .CK(debug_c_c), .Q(quadA_delayed[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(quadA_delayed[1]), .CK(debug_c_c), .Q(quadA_delayed_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n4156[3]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n4156[4]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n4156[5]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n4156[6]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n4156[7]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n4156[8]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n4156[9]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n4156[10]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n4156[11]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    CCU2D add_1649_33 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n26217), .S0(n4156[30]), 
          .S1(n4156[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1649_33.INIT0 = 16'h6969;
    defparam add_1649_33.INIT1 = 16'h6969;
    defparam add_1649_33.INJECT1_0 = "NO";
    defparam add_1649_33.INJECT1_1 = "NO";
    FD1P3IX count__i12 (.D(n4156[12]), .SP(n14013), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (debug_c_c, n8890, n32383, databus, 
            n608, n610, \control_reg[7] , n30314, Stepper_X_En_c, 
            Stepper_X_Dir_c, n13534, Stepper_X_M2_c_2, Stepper_X_M1_c_1, 
            \read_size[2] , n2644, n28137, n32384, n32381, n32382, 
            \read_size[0] , n21563, Stepper_X_M0_c_0, n579, prev_step_clk, 
            step_clk, prev_select, n30396, read_value, n9125, \register_addr[1] , 
            n11, \register_addr[0] , n30330, n3989, n30422, n30307, 
            n30489, n28421, n9118, limit_c_0, Stepper_X_Step_c, n34, 
            n26484, n24, n30313, n1, GND_net, VCC_net, Stepper_X_nFault_c, 
            n32380, n32385) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n8890;
    input n32383;
    input [31:0]databus;
    input n608;
    input n610;
    output \control_reg[7] ;
    input n30314;
    output Stepper_X_En_c;
    output Stepper_X_Dir_c;
    input n13534;
    output Stepper_X_M2_c_2;
    output Stepper_X_M1_c_1;
    output \read_size[2] ;
    input n2644;
    input n28137;
    input n32384;
    input n32381;
    input n32382;
    output \read_size[0] ;
    input n21563;
    output Stepper_X_M0_c_0;
    input n579;
    output prev_step_clk;
    output step_clk;
    output prev_select;
    input n30396;
    output [31:0]read_value;
    input n9125;
    input \register_addr[1] ;
    input n11;
    input \register_addr[0] ;
    output n30330;
    input n3989;
    input n30422;
    input n30307;
    input n30489;
    output n28421;
    output n9118;
    input limit_c_0;
    output Stepper_X_Step_c;
    input n34;
    output n26484;
    input n24;
    input n30313;
    input n1;
    input GND_net;
    input VCC_net;
    input Stepper_X_nFault_c;
    input n32380;
    input n32385;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n13511, n10750;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n3990;
    
    wire limit_latched, n182, prev_limit_latched, n41, n60, n54, 
        n42, n62, n28690, n52, n38, n58;
    wire [31:0]n100;
    
    wire n50_adj_27;
    wire [31:0]n224;
    
    wire n28691, n28692, n28693, int_step, n49, n56_adj_29, n46_adj_30, 
        n28631, n28632, n28633, n1_c, n2, n1_adj_31, n2_adj_32, 
        n1_adj_33, n2_adj_34, n1_adj_35, n2_adj_36, n2_adj_38, fault_latched, 
        n25966, n25965, n25964, n25963, n25962, n25961, n25960, 
        n25959, n25958, n25957, n25956, n25955, n25954, n25953, 
        n25952, n25951, n28688, n28689;
    
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n8890), .PD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n8890), .PD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n8890), .PD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n8890), .PD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n8890), .PD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n8890), .PD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n8890), .PD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n13511), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n13511), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n30314), .CD(n10750), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n30314), .PD(n32383), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n30314), .PD(n32383), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n13534), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n30314), .PD(n32383), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n13534), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n30314), .PD(n32383), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n28137), .SP(n2644), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3990[0]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3990[31]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3990[30]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3990[29]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n21563), .SP(n2644), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3990[28]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3990[27]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3990[26]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3990[25]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3990[24]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3990[23]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n13534), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13511), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n30396), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3990[22]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3990[21]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3990[20]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3990[19]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3990[18]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3990[17]), .CK(debug_c_c), .CD(n32383), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3990[16]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3990[15]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3990[14]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3990[13]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3990[12]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3990[11]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3990[10]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3990[9]), .CK(debug_c_c), .CD(n32384), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3990[8]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3990[7]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3990[6]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    FD1S3IX steps_reg__i5 (.D(n3990[5]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3990[4]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3990[3]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3990[2]), .CK(debug_c_c), .CD(n32381), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3990[1]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n28690), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i26_4_lut (.A(steps_reg[15]), .B(n52), .C(n38), .D(steps_reg[11]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_321 (.A(\register_addr[1] ), .B(n11), .C(\register_addr[0] ), 
         .Z(n30330)) /* synthesis lut_function=((B+(C))+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam i2_3_lut_rep_321.init = 16'hfdfd;
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    LUT4 i18_4_lut (.A(steps_reg[18]), .B(steps_reg[8]), .C(steps_reg[2]), 
         .D(steps_reg[16]), .Z(n50_adj_27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 mux_1589_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3989), .Z(n3990[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i1_3_lut.init = 16'hcaca;
    PFUMX i21540 (.BLUT(n28691), .ALUT(n28692), .C0(\register_addr[1] ), 
          .Z(n28693));
    LUT4 mux_1589_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3989), 
         .Z(n3990[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i32_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut (.A(n30422), .B(n30307), .C(n30489), .D(n28421), .Z(n9118)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0400;
    LUT4 mux_1589_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3989), 
         .Z(n3990[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3989), 
         .Z(n3990[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3989), 
         .Z(n3990[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3989), 
         .Z(n3990[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3989), 
         .Z(n3990[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3989), 
         .Z(n3990[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3989), 
         .Z(n3990[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3989), 
         .Z(n3990[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i24_3_lut.init = 16'hcaca;
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 mux_1589_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3989), 
         .Z(n3990[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3989), 
         .Z(n3990[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3989), 
         .Z(n3990[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3989), 
         .Z(n3990[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3989), 
         .Z(n3990[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3989), 
         .Z(n3990[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3989), 
         .Z(n3990[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3989), 
         .Z(n3990[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3989), 
         .Z(n3990[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3989), 
         .Z(n3990[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3989), 
         .Z(n3990[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3989), 
         .Z(n3990[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3989), 
         .Z(n3990[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3989), .Z(n3990[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3989), .Z(n3990[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3989), .Z(n3990[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3989), .Z(n3990[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3989), .Z(n3990[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3989), .Z(n3990[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3989), .Z(n3990[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3989), .Z(n3990[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1589_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3989), .Z(n3990[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1589_i2_3_lut.init = 16'hcaca;
    LUT4 i21274_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n28421)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21274_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i21538_3_lut (.A(Stepper_X_M2_c_2), .B(n34), .C(\register_addr[0] ), 
         .Z(n28691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21538_3_lut.init = 16'hcaca;
    LUT4 i21539_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n28692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21539_3_lut.init = 16'hcaca;
    LUT4 i9_2_lut (.A(steps_reg[24]), .B(steps_reg[1]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50_adj_27), .Z(n26484)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg[27]), .C(steps_reg[31]), 
         .D(steps_reg[30]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i28_4_lut (.A(steps_reg[6]), .B(n56_adj_29), .C(n46_adj_30), 
         .D(steps_reg[10]), .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[7]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[4]), .B(steps_reg[21]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[19]), .B(steps_reg[3]), .C(steps_reg[22]), 
         .D(steps_reg[13]), .Z(n56_adj_29)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[20]), .B(steps_reg[14]), .Z(n46_adj_30)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[29]), .B(steps_reg[12]), .C(steps_reg[9]), 
         .D(steps_reg[17]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    PFUMX i21480 (.BLUT(n28631), .ALUT(n28632), .C0(\register_addr[1] ), 
          .Z(n28633));
    LUT4 i6_2_lut (.A(steps_reg[28]), .B(steps_reg[23]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i15056_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15056_4_lut.init = 16'hc088;
    LUT4 i15057_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15057_4_lut.init = 16'hc088;
    PFUMX mux_1895_Mux_3_i3 (.BLUT(n1_c), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    LUT4 i15058_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15058_4_lut.init = 16'hc088;
    LUT4 i15059_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15059_4_lut.init = 16'hc088;
    PFUMX mux_1895_Mux_4_i3 (.BLUT(n1_adj_31), .ALUT(n2_adj_32), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    FD1P3AX int_step_182 (.D(n30313), .SP(n24), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i15060_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15060_4_lut.init = 16'hc088;
    PFUMX mux_1895_Mux_5_i3 (.BLUT(n1_adj_33), .ALUT(n2_adj_34), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    LUT4 i15061_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15061_4_lut.init = 16'hc088;
    PFUMX mux_1895_Mux_6_i3 (.BLUT(n1_adj_35), .ALUT(n2_adj_36), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    LUT4 i15062_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15062_4_lut.init = 16'hc088;
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    PFUMX mux_1895_Mux_7_i3 (.BLUT(n1), .ALUT(n2_adj_38), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    LUT4 i15063_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15063_4_lut.init = 16'hc088;
    LUT4 i15064_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15064_4_lut.init = 16'hc088;
    LUT4 i15065_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15065_4_lut.init = 16'hc088;
    LUT4 i15066_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15066_4_lut.init = 16'hc088;
    LUT4 i15067_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15067_4_lut.init = 16'hc088;
    LUT4 i15068_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15068_4_lut.init = 16'hc088;
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n28693), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n28633), .SP(n2644), .CD(n9125), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i15076_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15076_4_lut.init = 16'hc088;
    LUT4 i15077_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15077_4_lut.init = 16'hc088;
    LUT4 i15080_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15080_4_lut.init = 16'hc088;
    LUT4 i15081_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15081_4_lut.init = 16'hc088;
    LUT4 i15082_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15082_4_lut.init = 16'hc088;
    LUT4 i15083_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15083_4_lut.init = 16'hc088;
    LUT4 i15091_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15091_4_lut.init = 16'hc088;
    LUT4 i15092_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15092_4_lut.init = 16'hc088;
    LUT4 i21478_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n28631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21478_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25966), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25965), .COUT(n25966), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25964), .COUT(n25965), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25963), .COUT(n25964), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25962), .COUT(n25963), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25961), .COUT(n25962), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25960), .COUT(n25961), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25959), .COUT(n25960), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25958), .COUT(n25959), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25957), .COUT(n25958), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25956), .COUT(n25957), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25955), .COUT(n25956), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25954), .COUT(n25955), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25953), .COUT(n25954), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25952), .COUT(n25953), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25951), .COUT(n25952), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n34), .D1(prev_step_clk), 
          .COUT(n25951), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i21479_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n28632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21479_3_lut.init = 16'hcaca;
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    LUT4 i14870_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1_c)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14870_2_lut.init = 16'h2222;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    LUT4 mux_1895_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1895_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i14869_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_31)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14869_2_lut.init = 16'h2222;
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    LUT4 mux_1895_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2_adj_32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1895_Mux_4_i2_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n13511), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    LUT4 i14864_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_33)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14864_2_lut.init = 16'h2222;
    LUT4 mux_1895_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2_adj_34)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1895_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 i21535_3_lut (.A(Stepper_X_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n28688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21535_3_lut.init = 16'hcaca;
    LUT4 i14863_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_35)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14863_2_lut.init = 16'h2222;
    LUT4 mux_1895_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1895_Mux_6_i2_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n13511), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i15093_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15093_4_lut.init = 16'hc088;
    LUT4 i21536_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n28689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21536_3_lut.init = 16'hcaca;
    LUT4 mux_1895_Mux_7_i2_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), 
         .C(\register_addr[0] ), .Z(n2_adj_38)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1895_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_8 (.A(n8890), .B(n32380), .Z(n13511)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_8.init = 16'heeee;
    LUT4 i4343_3_lut (.A(prev_limit_latched), .B(n32380), .C(limit_latched), 
         .Z(n10750)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i4343_3_lut.init = 16'hdcdc;
    LUT4 i15094_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15094_4_lut.init = 16'hc088;
    LUT4 i15095_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15095_4_lut.init = 16'hc088;
    PFUMX i21537 (.BLUT(n28688), .ALUT(n28689), .C0(\register_addr[1] ), 
          .Z(n28690));
    ClockDivider_U8 step_clk_gen (.div_factor_reg({div_factor_reg}), .GND_net(GND_net), 
            .step_clk(step_clk), .debug_c_c(debug_c_c), .n32385(n32385), 
            .n32380(n32380)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (div_factor_reg, GND_net, step_clk, debug_c_c, 
            n32385, n32380) /* synthesis syn_module_defined=1 */ ;
    input [31:0]div_factor_reg;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n32385;
    input n32380;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25759, n25760, n25758, n25757, n25756, n25755, n25754, 
        n25753, n25752, n25751, n7643;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n30299;
    wire [31:0]n134;
    
    wire n25798, n7678, n25797;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n25796, n25795, n16283, n25794, n25793, n25792, n25791, 
        n25790, n25789, n25788, n25787, n25786, n25785, n26086, 
        n26085, n25784, n25783, n26084, n7712, n26083, n26082, 
        n25782;
    wire [31:0]n40;
    
    wire n26081, n26080, n26079, n26078, n26077, n25781, n25780, 
        n25779, n25778, n26076, n26075, n26074, n25777, n25776, 
        n26073, n26072, n26071, n25775, n25774, n25902, n25901, 
        n25900, n25899, n25773, n25772, n25898, n25897, n25771, 
        n25896, n25770, n25769, n25768, n25895, n25894, n25893, 
        n25767, n25892, n25766, n25891, n25890, n25765, n25889, 
        n25888, n25764, n25887, n25763, n25762, n25761;
    
    CCU2D sub_2017_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25759), .COUT(n25760));
    defparam sub_2017_add_2_19.INIT0 = 16'hf555;
    defparam sub_2017_add_2_19.INIT1 = 16'hf555;
    defparam sub_2017_add_2_19.INJECT1_0 = "NO";
    defparam sub_2017_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25758), .COUT(n25759));
    defparam sub_2017_add_2_17.INIT0 = 16'hf555;
    defparam sub_2017_add_2_17.INIT1 = 16'hf555;
    defparam sub_2017_add_2_17.INJECT1_0 = "NO";
    defparam sub_2017_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25757), .COUT(n25758));
    defparam sub_2017_add_2_15.INIT0 = 16'hf555;
    defparam sub_2017_add_2_15.INIT1 = 16'hf555;
    defparam sub_2017_add_2_15.INJECT1_0 = "NO";
    defparam sub_2017_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25756), .COUT(n25757));
    defparam sub_2017_add_2_13.INIT0 = 16'hf555;
    defparam sub_2017_add_2_13.INIT1 = 16'hf555;
    defparam sub_2017_add_2_13.INJECT1_0 = "NO";
    defparam sub_2017_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25755), .COUT(n25756));
    defparam sub_2017_add_2_11.INIT0 = 16'hf555;
    defparam sub_2017_add_2_11.INIT1 = 16'hf555;
    defparam sub_2017_add_2_11.INJECT1_0 = "NO";
    defparam sub_2017_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25754), .COUT(n25755));
    defparam sub_2017_add_2_9.INIT0 = 16'hf555;
    defparam sub_2017_add_2_9.INIT1 = 16'hf555;
    defparam sub_2017_add_2_9.INJECT1_0 = "NO";
    defparam sub_2017_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25753), .COUT(n25754));
    defparam sub_2017_add_2_7.INIT0 = 16'hf555;
    defparam sub_2017_add_2_7.INIT1 = 16'hf555;
    defparam sub_2017_add_2_7.INJECT1_0 = "NO";
    defparam sub_2017_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25752), .COUT(n25753));
    defparam sub_2017_add_2_5.INIT0 = 16'hf555;
    defparam sub_2017_add_2_5.INIT1 = 16'hf555;
    defparam sub_2017_add_2_5.INJECT1_0 = "NO";
    defparam sub_2017_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25751), .COUT(n25752));
    defparam sub_2017_add_2_3.INIT0 = 16'hf555;
    defparam sub_2017_add_2_3.INIT1 = 16'hf555;
    defparam sub_2017_add_2_3.INJECT1_0 = "NO";
    defparam sub_2017_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n25751));
    defparam sub_2017_add_2_1.INIT0 = 16'h0000;
    defparam sub_2017_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2017_add_2_1.INJECT1_0 = "NO";
    defparam sub_2017_add_2_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7643), .CK(debug_c_c), .CD(n32385), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2611__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i0.GSR = "ENABLED";
    CCU2D sub_2014_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25798), .S1(n7643));
    defparam sub_2014_add_2_33.INIT0 = 16'h5555;
    defparam sub_2014_add_2_33.INIT1 = 16'h0000;
    defparam sub_2014_add_2_33.INJECT1_0 = "NO";
    defparam sub_2014_add_2_33.INJECT1_1 = "NO";
    LUT4 i1009_2_lut_rep_290 (.A(n7678), .B(n32380), .Z(n30299)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1009_2_lut_rep_290.init = 16'heeee;
    CCU2D sub_2014_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25797), .COUT(n25798));
    defparam sub_2014_add_2_31.INIT0 = 16'h5999;
    defparam sub_2014_add_2_31.INIT1 = 16'h5999;
    defparam sub_2014_add_2_31.INJECT1_0 = "NO";
    defparam sub_2014_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25796), .COUT(n25797));
    defparam sub_2014_add_2_29.INIT0 = 16'h5999;
    defparam sub_2014_add_2_29.INIT1 = 16'h5999;
    defparam sub_2014_add_2_29.INJECT1_0 = "NO";
    defparam sub_2014_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25795), .COUT(n25796));
    defparam sub_2014_add_2_27.INIT0 = 16'h5999;
    defparam sub_2014_add_2_27.INIT1 = 16'h5999;
    defparam sub_2014_add_2_27.INJECT1_0 = "NO";
    defparam sub_2014_add_2_27.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    CCU2D sub_2014_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25794), .COUT(n25795));
    defparam sub_2014_add_2_25.INIT0 = 16'h5999;
    defparam sub_2014_add_2_25.INIT1 = 16'h5999;
    defparam sub_2014_add_2_25.INJECT1_0 = "NO";
    defparam sub_2014_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25793), .COUT(n25794));
    defparam sub_2014_add_2_23.INIT0 = 16'h5999;
    defparam sub_2014_add_2_23.INIT1 = 16'h5999;
    defparam sub_2014_add_2_23.INJECT1_0 = "NO";
    defparam sub_2014_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25792), .COUT(n25793));
    defparam sub_2014_add_2_21.INIT0 = 16'h5999;
    defparam sub_2014_add_2_21.INIT1 = 16'h5999;
    defparam sub_2014_add_2_21.INJECT1_0 = "NO";
    defparam sub_2014_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25791), .COUT(n25792));
    defparam sub_2014_add_2_19.INIT0 = 16'h5999;
    defparam sub_2014_add_2_19.INIT1 = 16'h5999;
    defparam sub_2014_add_2_19.INJECT1_0 = "NO";
    defparam sub_2014_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25790), .COUT(n25791));
    defparam sub_2014_add_2_17.INIT0 = 16'h5999;
    defparam sub_2014_add_2_17.INIT1 = 16'h5999;
    defparam sub_2014_add_2_17.INJECT1_0 = "NO";
    defparam sub_2014_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25789), .COUT(n25790));
    defparam sub_2014_add_2_15.INIT0 = 16'h5999;
    defparam sub_2014_add_2_15.INIT1 = 16'h5999;
    defparam sub_2014_add_2_15.INJECT1_0 = "NO";
    defparam sub_2014_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25788), .COUT(n25789));
    defparam sub_2014_add_2_13.INIT0 = 16'h5999;
    defparam sub_2014_add_2_13.INIT1 = 16'h5999;
    defparam sub_2014_add_2_13.INJECT1_0 = "NO";
    defparam sub_2014_add_2_13.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n30299), .CD(n16283), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n30299), .PD(n16283), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2014_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25787), .COUT(n25788));
    defparam sub_2014_add_2_11.INIT0 = 16'h5999;
    defparam sub_2014_add_2_11.INIT1 = 16'h5999;
    defparam sub_2014_add_2_11.INJECT1_0 = "NO";
    defparam sub_2014_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25786), .COUT(n25787));
    defparam sub_2014_add_2_9.INIT0 = 16'h5999;
    defparam sub_2014_add_2_9.INIT1 = 16'h5999;
    defparam sub_2014_add_2_9.INJECT1_0 = "NO";
    defparam sub_2014_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25785), .COUT(n25786));
    defparam sub_2014_add_2_7.INIT0 = 16'h5999;
    defparam sub_2014_add_2_7.INIT1 = 16'h5999;
    defparam sub_2014_add_2_7.INJECT1_0 = "NO";
    defparam sub_2014_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26086), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_33.INIT1 = 16'h0000;
    defparam count_2611_add_4_33.INJECT1_0 = "NO";
    defparam count_2611_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26085), .COUT(n26086), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_31.INJECT1_0 = "NO";
    defparam count_2611_add_4_31.INJECT1_1 = "NO";
    FD1S3IX count_2611__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i1.GSR = "ENABLED";
    CCU2D sub_2014_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25784), .COUT(n25785));
    defparam sub_2014_add_2_5.INIT0 = 16'h5999;
    defparam sub_2014_add_2_5.INIT1 = 16'h5999;
    defparam sub_2014_add_2_5.INJECT1_0 = "NO";
    defparam sub_2014_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25783), .COUT(n25784));
    defparam sub_2014_add_2_3.INIT0 = 16'h5999;
    defparam sub_2014_add_2_3.INIT1 = 16'h5999;
    defparam sub_2014_add_2_3.INJECT1_0 = "NO";
    defparam sub_2014_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26084), .COUT(n26085), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_29.INJECT1_0 = "NO";
    defparam count_2611_add_4_29.INJECT1_1 = "NO";
    FD1S3IX count_2611__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i2.GSR = "ENABLED";
    FD1S3IX count_2611__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i3.GSR = "ENABLED";
    FD1S3IX count_2611__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i4.GSR = "ENABLED";
    FD1S3IX count_2611__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i5.GSR = "ENABLED";
    FD1S3IX count_2611__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i6.GSR = "ENABLED";
    FD1S3IX count_2611__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i7.GSR = "ENABLED";
    FD1S3IX count_2611__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i8.GSR = "ENABLED";
    FD1S3IX count_2611__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i9.GSR = "ENABLED";
    FD1S3IX count_2611__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i10.GSR = "ENABLED";
    FD1S3IX count_2611__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i11.GSR = "ENABLED";
    FD1S3IX count_2611__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i12.GSR = "ENABLED";
    FD1S3IX count_2611__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i13.GSR = "ENABLED";
    FD1S3IX count_2611__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i14.GSR = "ENABLED";
    FD1S3IX count_2611__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i15.GSR = "ENABLED";
    FD1S3IX count_2611__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i16.GSR = "ENABLED";
    FD1S3IX count_2611__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i17.GSR = "ENABLED";
    FD1S3IX count_2611__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i18.GSR = "ENABLED";
    FD1S3IX count_2611__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i19.GSR = "ENABLED";
    FD1S3IX count_2611__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i20.GSR = "ENABLED";
    FD1S3IX count_2611__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i21.GSR = "ENABLED";
    FD1S3IX count_2611__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i22.GSR = "ENABLED";
    FD1S3IX count_2611__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i23.GSR = "ENABLED";
    FD1S3IX count_2611__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i24.GSR = "ENABLED";
    FD1S3IX count_2611__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i25.GSR = "ENABLED";
    FD1S3IX count_2611__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i26.GSR = "ENABLED";
    FD1S3IX count_2611__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i27.GSR = "ENABLED";
    FD1S3IX count_2611__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i28.GSR = "ENABLED";
    FD1S3IX count_2611__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i29.GSR = "ENABLED";
    FD1S3IX count_2611__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i30.GSR = "ENABLED";
    FD1S3IX count_2611__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n30299), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611__i31.GSR = "ENABLED";
    LUT4 i9900_2_lut_3_lut (.A(n7678), .B(n32380), .C(n7712), .Z(n16283)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9900_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_2014_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n25783));
    defparam sub_2014_add_2_1.INIT0 = 16'h0000;
    defparam sub_2014_add_2_1.INIT1 = 16'h5999;
    defparam sub_2014_add_2_1.INJECT1_0 = "NO";
    defparam sub_2014_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26083), .COUT(n26084), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_27.INJECT1_0 = "NO";
    defparam count_2611_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26082), .COUT(n26083), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_25.INJECT1_0 = "NO";
    defparam count_2611_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25782), .S1(n7678));
    defparam sub_2016_add_2_33.INIT0 = 16'h5999;
    defparam sub_2016_add_2_33.INIT1 = 16'h0000;
    defparam sub_2016_add_2_33.INJECT1_0 = "NO";
    defparam sub_2016_add_2_33.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26081), .COUT(n26082), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_23.INJECT1_0 = "NO";
    defparam count_2611_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26080), .COUT(n26081), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_21.INJECT1_0 = "NO";
    defparam count_2611_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26079), .COUT(n26080), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_19.INJECT1_0 = "NO";
    defparam count_2611_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26078), .COUT(n26079), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_17.INJECT1_0 = "NO";
    defparam count_2611_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26077), .COUT(n26078), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_15.INJECT1_0 = "NO";
    defparam count_2611_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25781), .COUT(n25782));
    defparam sub_2016_add_2_31.INIT0 = 16'h5999;
    defparam sub_2016_add_2_31.INIT1 = 16'h5999;
    defparam sub_2016_add_2_31.INJECT1_0 = "NO";
    defparam sub_2016_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25780), .COUT(n25781));
    defparam sub_2016_add_2_29.INIT0 = 16'h5999;
    defparam sub_2016_add_2_29.INIT1 = 16'h5999;
    defparam sub_2016_add_2_29.INJECT1_0 = "NO";
    defparam sub_2016_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25779), .COUT(n25780));
    defparam sub_2016_add_2_27.INIT0 = 16'h5999;
    defparam sub_2016_add_2_27.INIT1 = 16'h5999;
    defparam sub_2016_add_2_27.INJECT1_0 = "NO";
    defparam sub_2016_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25778), .COUT(n25779));
    defparam sub_2016_add_2_25.INIT0 = 16'h5999;
    defparam sub_2016_add_2_25.INIT1 = 16'h5999;
    defparam sub_2016_add_2_25.INJECT1_0 = "NO";
    defparam sub_2016_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26076), .COUT(n26077), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_13.INJECT1_0 = "NO";
    defparam count_2611_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26075), .COUT(n26076), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_11.INJECT1_0 = "NO";
    defparam count_2611_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26074), .COUT(n26075), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_9.INJECT1_0 = "NO";
    defparam count_2611_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25777), .COUT(n25778));
    defparam sub_2016_add_2_23.INIT0 = 16'h5999;
    defparam sub_2016_add_2_23.INIT1 = 16'h5999;
    defparam sub_2016_add_2_23.INJECT1_0 = "NO";
    defparam sub_2016_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25776), .COUT(n25777));
    defparam sub_2016_add_2_21.INIT0 = 16'h5999;
    defparam sub_2016_add_2_21.INIT1 = 16'h5999;
    defparam sub_2016_add_2_21.INJECT1_0 = "NO";
    defparam sub_2016_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26073), .COUT(n26074), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_7.INJECT1_0 = "NO";
    defparam count_2611_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26072), .COUT(n26073), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_5.INJECT1_0 = "NO";
    defparam count_2611_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26071), .COUT(n26072), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2611_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2611_add_4_3.INJECT1_0 = "NO";
    defparam count_2611_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2611_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26071), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2611_add_4_1.INIT0 = 16'hF000;
    defparam count_2611_add_4_1.INIT1 = 16'h0555;
    defparam count_2611_add_4_1.INJECT1_0 = "NO";
    defparam count_2611_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25775), .COUT(n25776));
    defparam sub_2016_add_2_19.INIT0 = 16'h5999;
    defparam sub_2016_add_2_19.INIT1 = 16'h5999;
    defparam sub_2016_add_2_19.INJECT1_0 = "NO";
    defparam sub_2016_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25774), .COUT(n25775));
    defparam sub_2016_add_2_17.INIT0 = 16'h5999;
    defparam sub_2016_add_2_17.INIT1 = 16'h5999;
    defparam sub_2016_add_2_17.INJECT1_0 = "NO";
    defparam sub_2016_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25902), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25901), .COUT(n25902), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25900), .COUT(n25901), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25899), .COUT(n25900), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25773), .COUT(n25774));
    defparam sub_2016_add_2_15.INIT0 = 16'h5999;
    defparam sub_2016_add_2_15.INIT1 = 16'h5999;
    defparam sub_2016_add_2_15.INJECT1_0 = "NO";
    defparam sub_2016_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25772), .COUT(n25773));
    defparam sub_2016_add_2_13.INIT0 = 16'h5999;
    defparam sub_2016_add_2_13.INIT1 = 16'h5999;
    defparam sub_2016_add_2_13.INJECT1_0 = "NO";
    defparam sub_2016_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25898), .COUT(n25899), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25897), .COUT(n25898), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25771), .COUT(n25772));
    defparam sub_2016_add_2_11.INIT0 = 16'h5999;
    defparam sub_2016_add_2_11.INIT1 = 16'h5999;
    defparam sub_2016_add_2_11.INJECT1_0 = "NO";
    defparam sub_2016_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25896), .COUT(n25897), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25770), .COUT(n25771));
    defparam sub_2016_add_2_9.INIT0 = 16'h5999;
    defparam sub_2016_add_2_9.INIT1 = 16'h5999;
    defparam sub_2016_add_2_9.INJECT1_0 = "NO";
    defparam sub_2016_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25769), .COUT(n25770));
    defparam sub_2016_add_2_7.INIT0 = 16'h5999;
    defparam sub_2016_add_2_7.INIT1 = 16'h5999;
    defparam sub_2016_add_2_7.INJECT1_0 = "NO";
    defparam sub_2016_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25768), .COUT(n25769));
    defparam sub_2016_add_2_5.INIT0 = 16'h5999;
    defparam sub_2016_add_2_5.INIT1 = 16'h5999;
    defparam sub_2016_add_2_5.INJECT1_0 = "NO";
    defparam sub_2016_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25895), .COUT(n25896), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25894), .COUT(n25895), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25893), .COUT(n25894), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25767), .COUT(n25768));
    defparam sub_2016_add_2_3.INIT0 = 16'h5999;
    defparam sub_2016_add_2_3.INIT1 = 16'h5999;
    defparam sub_2016_add_2_3.INJECT1_0 = "NO";
    defparam sub_2016_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n25767));
    defparam sub_2016_add_2_1.INIT0 = 16'h0000;
    defparam sub_2016_add_2_1.INIT1 = 16'h5999;
    defparam sub_2016_add_2_1.INJECT1_0 = "NO";
    defparam sub_2016_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25892), .COUT(n25893), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25766), .S1(n7712));
    defparam sub_2017_add_2_33.INIT0 = 16'hf555;
    defparam sub_2017_add_2_33.INIT1 = 16'h0000;
    defparam sub_2017_add_2_33.INJECT1_0 = "NO";
    defparam sub_2017_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25891), .COUT(n25892), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25890), .COUT(n25891), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25765), .COUT(n25766));
    defparam sub_2017_add_2_31.INIT0 = 16'hf555;
    defparam sub_2017_add_2_31.INIT1 = 16'hf555;
    defparam sub_2017_add_2_31.INJECT1_0 = "NO";
    defparam sub_2017_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25889), .COUT(n25890), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25888), .COUT(n25889), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25764), .COUT(n25765));
    defparam sub_2017_add_2_29.INIT0 = 16'hf555;
    defparam sub_2017_add_2_29.INIT1 = 16'hf555;
    defparam sub_2017_add_2_29.INJECT1_0 = "NO";
    defparam sub_2017_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25887), .COUT(n25888), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25887), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25763), .COUT(n25764));
    defparam sub_2017_add_2_27.INIT0 = 16'hf555;
    defparam sub_2017_add_2_27.INIT1 = 16'hf555;
    defparam sub_2017_add_2_27.INJECT1_0 = "NO";
    defparam sub_2017_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25762), .COUT(n25763));
    defparam sub_2017_add_2_25.INIT0 = 16'hf555;
    defparam sub_2017_add_2_25.INIT1 = 16'hf555;
    defparam sub_2017_add_2_25.INJECT1_0 = "NO";
    defparam sub_2017_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25761), .COUT(n25762));
    defparam sub_2017_add_2_23.INIT0 = 16'hf555;
    defparam sub_2017_add_2_23.INIT1 = 16'hf555;
    defparam sub_2017_add_2_23.INJECT1_0 = "NO";
    defparam sub_2017_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2017_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25760), .COUT(n25761));
    defparam sub_2017_add_2_21.INIT0 = 16'hf555;
    defparam sub_2017_add_2_21.INIT1 = 16'hf555;
    defparam sub_2017_add_2_21.INJECT1_0 = "NO";
    defparam sub_2017_add_2_21.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (read_value, debug_c_c, n2673, 
            n9136, n32382, VCC_net, GND_net, Stepper_A_nFault_c, \read_size[0] , 
            n28324, Stepper_A_M0_c_0, databus, prev_select, n30371, 
            n32383, n32381, \control_reg[7] , Stepper_A_En_c, Stepper_A_Dir_c, 
            Stepper_A_M2_c_2, Stepper_A_M1_c_1, \register_addr[0] , n3806, 
            \register_addr[1] , stepping, n26585, \steps_reg[7] , \register_addr[5] , 
            \register_addr[4] , n21533, limit_c_3, Stepper_A_Step_c, 
            n30491, n28218, rw, n30338, n13269, n28184, n30411, 
            n32380, \read_size[2] , n28172, n32, prev_step_clk, step_clk, 
            n30310, n32385, n32386, n22, n32_adj_1, prev_step_clk_adj_2, 
            step_clk_adj_3, n30311, n22_adj_4, prev_step_clk_adj_5, 
            n34, step_clk_adj_6, n30313, n24, n19) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2673;
    input n9136;
    input n32382;
    input VCC_net;
    input GND_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n28324;
    output Stepper_A_M0_c_0;
    input [31:0]databus;
    output prev_select;
    input n30371;
    input n32383;
    input n32381;
    output \control_reg[7] ;
    output Stepper_A_En_c;
    output Stepper_A_Dir_c;
    output Stepper_A_M2_c_2;
    output Stepper_A_M1_c_1;
    input \register_addr[0] ;
    input n3806;
    input \register_addr[1] ;
    input stepping;
    output n26585;
    output \steps_reg[7] ;
    input \register_addr[5] ;
    input \register_addr[4] ;
    output n21533;
    input limit_c_3;
    output Stepper_A_Step_c;
    input n30491;
    output n28218;
    input rw;
    input n30338;
    input n13269;
    input n28184;
    input n30411;
    input n32380;
    output \read_size[2] ;
    input n28172;
    input n32;
    input prev_step_clk;
    input step_clk;
    output n30310;
    input n32385;
    input n32386;
    output n22;
    input n32_adj_1;
    input prev_step_clk_adj_2;
    input step_clk_adj_3;
    output n30311;
    output n22_adj_4;
    input prev_step_clk_adj_5;
    input n34;
    input step_clk_adj_6;
    output n30313;
    output n24;
    input n19;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n28678;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n3807;
    
    wire fault_latched, n13605, prev_step_clk_c, step_clk_c, limit_latched, 
        n182, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n8919, n11663;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n28646, n28647, n28648;
    wire [31:0]n100;
    
    wire n18628, n28681;
    wire [31:0]n224;
    
    wire n49, n62_adj_1, n58_adj_2, n50_adj_3, n41, n60_adj_4, n54_adj_5, 
        n42_adj_6, n52_adj_7, n38_adj_8, n56_adj_9, n46_adj_10, int_step, 
        n28676, n28677, n13, n30312, n30;
    wire [31:0]n99;
    
    wire n18626, n28679, n28680, n25918, n25917, n25916, n25915, 
        n25914, n25913, n25912, n25911, n25910, n25909, n25908, 
        n25907, n25906, n25905, n25904, n25903;
    wire [7:0]n8280;
    wire [31:0]n7169;
    
    FD1P3IX read_value__i0 (.D(n28678), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3807[0]), .CK(debug_c_c), .CD(n32382), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n28324), .SP(n2673), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n13605), .CD(n32382), 
            .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk_c), .CK(debug_c_c), .Q(prev_step_clk_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n30371), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n8919), .CD(n32383), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n8919), .PD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n8919), .PD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n8919), .PD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n8919), .PD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n8919), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n8919), .PD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n8919), .PD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n8919), .PD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n8919), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n8919), .CD(n32381), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n8919), .CD(n32382), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13605), .CD(n11663), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13605), .PD(n32382), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13605), .PD(n32382), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13605), .CD(n32381), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13605), .PD(n32381), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13605), .CD(n32382), 
            .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13605), .PD(n32381), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    PFUMX i21495 (.BLUT(n28646), .ALUT(n28647), .C0(\register_addr[0] ), 
          .Z(n28648));
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n18628), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n28648), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n28681), .SP(n2673), .CD(n9136), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1542_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3806), 
         .Z(n3807[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3806), 
         .Z(n3807[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3806), 
         .Z(n3807[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3806), .Z(n3807[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3806), 
         .Z(n3807[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3806), 
         .Z(n3807[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i28_3_lut.init = 16'hcaca;
    LUT4 i21493_3_lut (.A(Stepper_A_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n28646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21493_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3806), 
         .Z(n3807[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i27_3_lut.init = 16'hcaca;
    LUT4 i21494_3_lut (.A(stepping), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n28647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21494_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3806), 
         .Z(n3807[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3806), 
         .Z(n3807[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3806), 
         .Z(n3807[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3806), 
         .Z(n3807[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3806), 
         .Z(n3807[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3806), 
         .Z(n3807[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3806), 
         .Z(n3807[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3806), 
         .Z(n3807[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3806), 
         .Z(n3807[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3806), 
         .Z(n3807[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i17_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_1), .C(n58_adj_2), .D(n50_adj_3), 
         .Z(n26585)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[18]), .B(steps_reg[12]), .C(steps_reg[28]), 
         .D(steps_reg[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 mux_1542_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3806), 
         .Z(n3807[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i16_3_lut.init = 16'hcaca;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_4), .C(n54_adj_5), .D(n42_adj_6), 
         .Z(n62_adj_1)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 mux_1542_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3806), 
         .Z(n3807[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i15_3_lut.init = 16'hcaca;
    LUT4 i26_4_lut (.A(steps_reg[9]), .B(n52_adj_7), .C(n38_adj_8), .D(steps_reg[27]), 
         .Z(n58_adj_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 mux_1542_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3806), 
         .Z(n3807[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i14_3_lut.init = 16'hcaca;
    LUT4 i18_4_lut (.A(steps_reg[11]), .B(steps_reg[25]), .C(steps_reg[21]), 
         .D(steps_reg[26]), .Z(n50_adj_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 mux_1542_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3806), 
         .Z(n3807[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3806), 
         .Z(n3807[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3806), 
         .Z(n3807[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i11_3_lut.init = 16'hcaca;
    LUT4 i9_2_lut (.A(steps_reg[5]), .B(steps_reg[15]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[3]), .B(n56_adj_9), .C(n46_adj_10), .D(steps_reg[31]), 
         .Z(n60_adj_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 mux_1542_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3806), .Z(n3807[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3806), .Z(n3807[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3806), .Z(n3807[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i8_3_lut.init = 16'hcaca;
    LUT4 i22_4_lut (.A(steps_reg[13]), .B(steps_reg[0]), .C(steps_reg[17]), 
         .D(steps_reg[24]), .Z(n54_adj_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 mux_1542_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3806), .Z(n3807[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i7_3_lut.init = 16'hcaca;
    LUT4 i10_2_lut (.A(steps_reg[23]), .B(steps_reg[29]), .Z(n42_adj_6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[8]), .B(steps_reg[2]), .C(steps_reg[16]), 
         .D(steps_reg[4]), .Z(n56_adj_9)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[6]), .B(steps_reg[20]), .Z(n46_adj_10)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 mux_1542_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3806), .Z(n3807[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i6_3_lut.init = 16'hcaca;
    LUT4 i20_4_lut (.A(steps_reg[14]), .B(steps_reg[22]), .C(steps_reg[19]), 
         .D(steps_reg[1]), .Z(n52_adj_7)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 mux_1542_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3806), .Z(n3807[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3806), .Z(n3807[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3806), .Z(n3807[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3806), .Z(n3807[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1542_i2_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut (.A(steps_reg[30]), .B(\steps_reg[7] ), .Z(n38_adj_8)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i15155_2_lut (.A(\register_addr[5] ), .B(\register_addr[4] ), .Z(n21533)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15155_2_lut.init = 16'h8888;
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i21523_3_lut (.A(Stepper_A_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n28676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21523_3_lut.init = 16'hcaca;
    LUT4 i21524_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n28677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21524_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(n30491), .D(\register_addr[4] ), .Z(n28218)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0002;
    LUT4 i21681_2_lut_3_lut_4_lut (.A(rw), .B(n30338), .C(n21533), .D(n13269), 
         .Z(n13605)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i21681_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i2_3_lut_4_lut (.A(rw), .B(n30338), .C(n28184), .D(n30411), 
         .Z(n8919)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_4_lut.init = 16'h4000;
    LUT4 i5256_3_lut (.A(prev_limit_latched), .B(n32380), .C(limit_latched), 
         .Z(n11663)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i5256_3_lut.init = 16'hdcdc;
    FD1P3AX int_step_182 (.D(n30312), .SP(n13), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n28172), .SP(n2673), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_301 (.A(n32), .B(prev_step_clk), .C(step_clk), .Z(n30310)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_301.init = 16'h2020;
    LUT4 i1_4_lut (.A(div_factor_reg[10]), .B(n30), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n99[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_adj_1 (.A(\register_addr[1] ), .B(n9136), .Z(n30)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_2_lut_adj_1.init = 16'h2222;
    LUT4 i1_4_lut_adj_2 (.A(div_factor_reg[11]), .B(n30), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n99[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_2.init = 16'hc088;
    LUT4 i1_4_lut_adj_3 (.A(div_factor_reg[12]), .B(n30), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n99[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_3.init = 16'hc088;
    FD1S3IX steps_reg__i31 (.D(n3807[31]), .CK(debug_c_c), .CD(n32385), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3807[30]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3807[29]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3807[28]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3807[27]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3807[26]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3807[25]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3807[24]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3807[23]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3807[22]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3807[21]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3807[20]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3807[19]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3807[18]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3807[17]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3807[16]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3807[15]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3807[14]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3807[13]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3807[12]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3807[11]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3807[10]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3807[9]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3807[8]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3807[7]), .CK(debug_c_c), .CD(n32386), 
            .Q(\steps_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3807[6]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3807[5]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3807[4]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3807[3]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3807[2]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3807[1]), .CK(debug_c_c), .CD(n32386), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i14595_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14595_4_lut.init = 16'hc088;
    LUT4 i14596_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14596_4_lut.init = 16'hc088;
    LUT4 i14597_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14597_4_lut.init = 16'hc088;
    LUT4 i14598_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14598_4_lut.init = 16'hc088;
    LUT4 i14599_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14599_4_lut.init = 16'hc088;
    LUT4 i14600_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14600_4_lut.init = 16'hc088;
    LUT4 i14601_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14601_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_4 (.A(\register_addr[1] ), .B(div_factor_reg[24]), 
         .C(steps_reg[24]), .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_4.init = 16'ha088;
    LUT4 i14602_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14602_4_lut.init = 16'hc088;
    LUT4 i14603_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14603_4_lut.init = 16'hc088;
    LUT4 i14604_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14604_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_5 (.A(\register_addr[1] ), .B(div_factor_reg[20]), 
         .C(steps_reg[20]), .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_5.init = 16'ha088;
    LUT4 i14605_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14605_4_lut.init = 16'hc088;
    LUT4 i14606_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14606_4_lut.init = 16'hc088;
    LUT4 i14607_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14607_4_lut.init = 16'hc088;
    LUT4 i14608_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14608_4_lut.init = 16'hc088;
    LUT4 i14609_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14609_4_lut.init = 16'hc088;
    LUT4 i14610_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14610_4_lut.init = 16'hc088;
    LUT4 i14611_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14611_4_lut.init = 16'hc088;
    LUT4 i14612_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14612_4_lut.init = 16'hc088;
    LUT4 i14613_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14613_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_4_lut (.A(n32), .B(prev_step_clk), .C(step_clk), .D(n32380), 
         .Z(n22)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut.init = 16'h002c;
    PFUMX i21525 (.BLUT(n28676), .ALUT(n28677), .C0(\register_addr[1] ), 
          .Z(n28678));
    LUT4 i2_3_lut_rep_302 (.A(n32_adj_1), .B(prev_step_clk_adj_2), .C(step_clk_adj_3), 
         .Z(n30311)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_302.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_adj_6 (.A(n32_adj_1), .B(prev_step_clk_adj_2), .C(step_clk_adj_3), 
         .D(n32380), .Z(n22_adj_4)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_6.init = 16'h002c;
    LUT4 i2_3_lut_rep_304 (.A(prev_step_clk_adj_5), .B(n34), .C(step_clk_adj_6), 
         .Z(n30313)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_304.init = 16'h4040;
    LUT4 i1_4_lut_4_lut_adj_7 (.A(prev_step_clk_adj_5), .B(n34), .C(step_clk_adj_6), 
         .D(n32380), .Z(n24)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_7.init = 16'h004a;
    FD1P3AX read_value__i10 (.D(n99[10]), .SP(n2673), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n99[11]), .SP(n2673), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n99[12]), .SP(n2673), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    LUT4 i12222_3_lut (.A(\control_reg[7] ), .B(div_factor_reg[7]), .C(\register_addr[1] ), 
         .Z(n18626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i12222_3_lut.init = 16'hcaca;
    LUT4 i21526_3_lut (.A(Stepper_A_M1_c_1), .B(div_factor_reg[1]), .C(\register_addr[1] ), 
         .Z(n28679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21526_3_lut.init = 16'hcaca;
    LUT4 i21527_3_lut (.A(fault_latched), .B(steps_reg[1]), .C(\register_addr[1] ), 
         .Z(n28680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21527_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25918), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25917), .COUT(n25918), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25916), .COUT(n25917), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25915), .COUT(n25916), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25914), .COUT(n25915), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25913), .COUT(n25914), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25912), .COUT(n25913), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25911), .COUT(n25912), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25910), .COUT(n25911), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25909), .COUT(n25910), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25908), .COUT(n25909), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25907), .COUT(n25908), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(\steps_reg[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25906), .COUT(n25907), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25905), .COUT(n25906), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    PFUMX i12224 (.BLUT(n18626), .ALUT(n19), .C0(\register_addr[0] ), 
          .Z(n18628));
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25904), .COUT(n25905), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25903), .COUT(n25904), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk_c), .C1(stepping), .D1(prev_step_clk_c), 
          .COUT(n25903), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    PFUMX i21528 (.BLUT(n28679), .ALUT(n28680), .C0(\register_addr[0] ), 
          .Z(n28681));
    LUT4 i14594_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8280[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14594_2_lut.init = 16'h2222;
    LUT4 mux_1967_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7169[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1967_i4_3_lut.init = 16'hcaca;
    LUT4 i14593_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8280[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14593_2_lut.init = 16'h2222;
    LUT4 mux_1967_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7169[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1967_i5_3_lut.init = 16'hcaca;
    LUT4 i14592_2_lut (.A(Stepper_A_Dir_c), .B(\register_addr[0] ), .Z(n8280[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14592_2_lut.init = 16'h2222;
    LUT4 mux_1967_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7169[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1967_i6_3_lut.init = 16'hcaca;
    LUT4 i14591_2_lut (.A(Stepper_A_En_c), .B(\register_addr[0] ), .Z(n8280[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14591_2_lut.init = 16'h2222;
    LUT4 mux_1967_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7169[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1967_i7_3_lut.init = 16'hcaca;
    PFUMX mux_1971_i4 (.BLUT(n8280[3]), .ALUT(n7169[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_1971_i5 (.BLUT(n8280[4]), .ALUT(n7169[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1971_i6 (.BLUT(n8280[5]), .ALUT(n7169[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1971_i7 (.BLUT(n8280[6]), .ALUT(n7169[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    ClockDivider_U9 step_clk_gen (.div_factor_reg({div_factor_reg}), .GND_net(GND_net), 
            .step_clk(step_clk_c), .debug_c_c(debug_c_c), .n32385(n32385), 
            .stepping(stepping), .prev_step_clk(prev_step_clk_c), .n30312(n30312), 
            .n32380(n32380), .n13(n13)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (div_factor_reg, GND_net, step_clk, debug_c_c, 
            n32385, stepping, prev_step_clk, n30312, n32380, n13) /* synthesis syn_module_defined=1 */ ;
    input [31:0]div_factor_reg;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n32385;
    input stepping;
    input prev_step_clk;
    output n30312;
    input n32380;
    output n13;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25607, n25608, n26047;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n26048, n26046, n26045, n26044, n26043, n26042, n26041, 
        n26040, n26039, n25654, n7955, n25653;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n25652, n25651, n25650, n25649, n25648, n25647, n30300, 
        n25646, n25645, n25854;
    wire [31:0]n40;
    
    wire n25853, n25852, n25851, n25850, n25849, n25848, n25847, 
        n25846, n25845, n25844, n25843, n25842, n25841, n25840, 
        n25839, n25644, n25643, n25642, n25641, n25640, n25639, 
        n25638, n7990, n25637, n25636, n25635, n25634, n25633, 
        n25632, n25631, n25630, n25629, n25628, n25627, n25626, 
        n25625, n25624, n25623, n25622, n8024, n25621, n16223, 
        n25620, n25619, n25618, n25617, n25616, n25615, n25614, 
        n25613, n25612, n26054, n26053, n25611, n26052, n26051, 
        n25610, n25609, n26050, n26049;
    
    CCU2D sub_2032_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25607), .COUT(n25608));
    defparam sub_2032_add_2_3.INIT0 = 16'hf555;
    defparam sub_2032_add_2_3.INIT1 = 16'hf555;
    defparam sub_2032_add_2_3.INJECT1_0 = "NO";
    defparam sub_2032_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26047), .COUT(n26048), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_19.INJECT1_0 = "NO";
    defparam count_2614_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26046), .COUT(n26047), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_17.INJECT1_0 = "NO";
    defparam count_2614_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26045), .COUT(n26046), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_15.INJECT1_0 = "NO";
    defparam count_2614_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26044), .COUT(n26045), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_13.INJECT1_0 = "NO";
    defparam count_2614_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26043), .COUT(n26044), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_11.INJECT1_0 = "NO";
    defparam count_2614_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26042), .COUT(n26043), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_9.INJECT1_0 = "NO";
    defparam count_2614_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26041), .COUT(n26042), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_7.INJECT1_0 = "NO";
    defparam count_2614_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n25607));
    defparam sub_2032_add_2_1.INIT0 = 16'h0000;
    defparam sub_2032_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2032_add_2_1.INJECT1_0 = "NO";
    defparam sub_2032_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26040), .COUT(n26041), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_5.INJECT1_0 = "NO";
    defparam count_2614_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26039), .COUT(n26040), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_3.INJECT1_0 = "NO";
    defparam count_2614_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26039), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_1.INIT0 = 16'hF000;
    defparam count_2614_add_4_1.INIT1 = 16'h0555;
    defparam count_2614_add_4_1.INJECT1_0 = "NO";
    defparam count_2614_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25654), .S1(n7955));
    defparam sub_2029_add_2_33.INIT0 = 16'h5555;
    defparam sub_2029_add_2_33.INIT1 = 16'h0000;
    defparam sub_2029_add_2_33.INJECT1_0 = "NO";
    defparam sub_2029_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25653), .COUT(n25654));
    defparam sub_2029_add_2_31.INIT0 = 16'h5999;
    defparam sub_2029_add_2_31.INIT1 = 16'h5999;
    defparam sub_2029_add_2_31.INJECT1_0 = "NO";
    defparam sub_2029_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25652), .COUT(n25653));
    defparam sub_2029_add_2_29.INIT0 = 16'h5999;
    defparam sub_2029_add_2_29.INIT1 = 16'h5999;
    defparam sub_2029_add_2_29.INJECT1_0 = "NO";
    defparam sub_2029_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25651), .COUT(n25652));
    defparam sub_2029_add_2_27.INIT0 = 16'h5999;
    defparam sub_2029_add_2_27.INIT1 = 16'h5999;
    defparam sub_2029_add_2_27.INJECT1_0 = "NO";
    defparam sub_2029_add_2_27.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7955), .CK(debug_c_c), .CD(n32385), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2029_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25650), .COUT(n25651));
    defparam sub_2029_add_2_25.INIT0 = 16'h5999;
    defparam sub_2029_add_2_25.INIT1 = 16'h5999;
    defparam sub_2029_add_2_25.INJECT1_0 = "NO";
    defparam sub_2029_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25649), .COUT(n25650));
    defparam sub_2029_add_2_23.INIT0 = 16'h5999;
    defparam sub_2029_add_2_23.INIT1 = 16'h5999;
    defparam sub_2029_add_2_23.INJECT1_0 = "NO";
    defparam sub_2029_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25648), .COUT(n25649));
    defparam sub_2029_add_2_21.INIT0 = 16'h5999;
    defparam sub_2029_add_2_21.INIT1 = 16'h5999;
    defparam sub_2029_add_2_21.INJECT1_0 = "NO";
    defparam sub_2029_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25647), .COUT(n25648));
    defparam sub_2029_add_2_19.INIT0 = 16'h5999;
    defparam sub_2029_add_2_19.INIT1 = 16'h5999;
    defparam sub_2029_add_2_19.INJECT1_0 = "NO";
    defparam sub_2029_add_2_19.INJECT1_1 = "NO";
    FD1S3IX count_2614__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i0.GSR = "ENABLED";
    CCU2D sub_2029_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25646), .COUT(n25647));
    defparam sub_2029_add_2_17.INIT0 = 16'h5999;
    defparam sub_2029_add_2_17.INIT1 = 16'h5999;
    defparam sub_2029_add_2_17.INJECT1_0 = "NO";
    defparam sub_2029_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25645), .COUT(n25646));
    defparam sub_2029_add_2_15.INIT0 = 16'h5999;
    defparam sub_2029_add_2_15.INIT1 = 16'h5999;
    defparam sub_2029_add_2_15.INJECT1_0 = "NO";
    defparam sub_2029_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25854), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25853), .COUT(n25854), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25852), .COUT(n25853), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25851), .COUT(n25852), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25850), .COUT(n25851), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25849), .COUT(n25850), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25848), .COUT(n25849), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25847), .COUT(n25848), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25846), .COUT(n25847), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25845), .COUT(n25846), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25844), .COUT(n25845), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25843), .COUT(n25844), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25842), .COUT(n25843), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25841), .COUT(n25842), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25840), .COUT(n25841), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25839), .COUT(n25840), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25839), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25644), .COUT(n25645));
    defparam sub_2029_add_2_13.INIT0 = 16'h5999;
    defparam sub_2029_add_2_13.INIT1 = 16'h5999;
    defparam sub_2029_add_2_13.INJECT1_0 = "NO";
    defparam sub_2029_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25643), .COUT(n25644));
    defparam sub_2029_add_2_11.INIT0 = 16'h5999;
    defparam sub_2029_add_2_11.INIT1 = 16'h5999;
    defparam sub_2029_add_2_11.INJECT1_0 = "NO";
    defparam sub_2029_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25642), .COUT(n25643));
    defparam sub_2029_add_2_9.INIT0 = 16'h5999;
    defparam sub_2029_add_2_9.INIT1 = 16'h5999;
    defparam sub_2029_add_2_9.INJECT1_0 = "NO";
    defparam sub_2029_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25641), .COUT(n25642));
    defparam sub_2029_add_2_7.INIT0 = 16'h5999;
    defparam sub_2029_add_2_7.INIT1 = 16'h5999;
    defparam sub_2029_add_2_7.INJECT1_0 = "NO";
    defparam sub_2029_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25640), .COUT(n25641));
    defparam sub_2029_add_2_5.INIT0 = 16'h5999;
    defparam sub_2029_add_2_5.INIT1 = 16'h5999;
    defparam sub_2029_add_2_5.INJECT1_0 = "NO";
    defparam sub_2029_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25639), .COUT(n25640));
    defparam sub_2029_add_2_3.INIT0 = 16'h5999;
    defparam sub_2029_add_2_3.INIT1 = 16'h5999;
    defparam sub_2029_add_2_3.INJECT1_0 = "NO";
    defparam sub_2029_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n25639));
    defparam sub_2029_add_2_1.INIT0 = 16'h0000;
    defparam sub_2029_add_2_1.INIT1 = 16'h5999;
    defparam sub_2029_add_2_1.INJECT1_0 = "NO";
    defparam sub_2029_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25638), .S1(n7990));
    defparam sub_2031_add_2_33.INIT0 = 16'h5999;
    defparam sub_2031_add_2_33.INIT1 = 16'h0000;
    defparam sub_2031_add_2_33.INJECT1_0 = "NO";
    defparam sub_2031_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25637), .COUT(n25638));
    defparam sub_2031_add_2_31.INIT0 = 16'h5999;
    defparam sub_2031_add_2_31.INIT1 = 16'h5999;
    defparam sub_2031_add_2_31.INJECT1_0 = "NO";
    defparam sub_2031_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25636), .COUT(n25637));
    defparam sub_2031_add_2_29.INIT0 = 16'h5999;
    defparam sub_2031_add_2_29.INIT1 = 16'h5999;
    defparam sub_2031_add_2_29.INJECT1_0 = "NO";
    defparam sub_2031_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25635), .COUT(n25636));
    defparam sub_2031_add_2_27.INIT0 = 16'h5999;
    defparam sub_2031_add_2_27.INIT1 = 16'h5999;
    defparam sub_2031_add_2_27.INJECT1_0 = "NO";
    defparam sub_2031_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25634), .COUT(n25635));
    defparam sub_2031_add_2_25.INIT0 = 16'h5999;
    defparam sub_2031_add_2_25.INIT1 = 16'h5999;
    defparam sub_2031_add_2_25.INJECT1_0 = "NO";
    defparam sub_2031_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25633), .COUT(n25634));
    defparam sub_2031_add_2_23.INIT0 = 16'h5999;
    defparam sub_2031_add_2_23.INIT1 = 16'h5999;
    defparam sub_2031_add_2_23.INJECT1_0 = "NO";
    defparam sub_2031_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25632), .COUT(n25633));
    defparam sub_2031_add_2_21.INIT0 = 16'h5999;
    defparam sub_2031_add_2_21.INIT1 = 16'h5999;
    defparam sub_2031_add_2_21.INJECT1_0 = "NO";
    defparam sub_2031_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25631), .COUT(n25632));
    defparam sub_2031_add_2_19.INIT0 = 16'h5999;
    defparam sub_2031_add_2_19.INIT1 = 16'h5999;
    defparam sub_2031_add_2_19.INJECT1_0 = "NO";
    defparam sub_2031_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25630), .COUT(n25631));
    defparam sub_2031_add_2_17.INIT0 = 16'h5999;
    defparam sub_2031_add_2_17.INIT1 = 16'h5999;
    defparam sub_2031_add_2_17.INJECT1_0 = "NO";
    defparam sub_2031_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25629), .COUT(n25630));
    defparam sub_2031_add_2_15.INIT0 = 16'h5999;
    defparam sub_2031_add_2_15.INIT1 = 16'h5999;
    defparam sub_2031_add_2_15.INJECT1_0 = "NO";
    defparam sub_2031_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25628), .COUT(n25629));
    defparam sub_2031_add_2_13.INIT0 = 16'h5999;
    defparam sub_2031_add_2_13.INIT1 = 16'h5999;
    defparam sub_2031_add_2_13.INJECT1_0 = "NO";
    defparam sub_2031_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n25627), .COUT(n25628));
    defparam sub_2031_add_2_11.INIT0 = 16'h5999;
    defparam sub_2031_add_2_11.INIT1 = 16'h5999;
    defparam sub_2031_add_2_11.INJECT1_0 = "NO";
    defparam sub_2031_add_2_11.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_303 (.A(stepping), .B(prev_step_clk), .C(step_clk), 
         .Z(n30312)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i2_3_lut_rep_303.init = 16'h2020;
    LUT4 i1_4_lut_4_lut (.A(stepping), .B(prev_step_clk), .C(step_clk), 
         .D(n32380), .Z(n13)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i1_4_lut_4_lut.init = 16'h002c;
    CCU2D sub_2031_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25626), .COUT(n25627));
    defparam sub_2031_add_2_9.INIT0 = 16'h5999;
    defparam sub_2031_add_2_9.INIT1 = 16'h5999;
    defparam sub_2031_add_2_9.INJECT1_0 = "NO";
    defparam sub_2031_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25625), .COUT(n25626));
    defparam sub_2031_add_2_7.INIT0 = 16'h5999;
    defparam sub_2031_add_2_7.INIT1 = 16'h5999;
    defparam sub_2031_add_2_7.INJECT1_0 = "NO";
    defparam sub_2031_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25624), .COUT(n25625));
    defparam sub_2031_add_2_5.INIT0 = 16'h5999;
    defparam sub_2031_add_2_5.INIT1 = 16'h5999;
    defparam sub_2031_add_2_5.INJECT1_0 = "NO";
    defparam sub_2031_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n25623), .COUT(n25624));
    defparam sub_2031_add_2_3.INIT0 = 16'h5999;
    defparam sub_2031_add_2_3.INIT1 = 16'h5999;
    defparam sub_2031_add_2_3.INJECT1_0 = "NO";
    defparam sub_2031_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2031_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n25623));
    defparam sub_2031_add_2_1.INIT0 = 16'h0000;
    defparam sub_2031_add_2_1.INIT1 = 16'h5999;
    defparam sub_2031_add_2_1.INJECT1_0 = "NO";
    defparam sub_2031_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25622), .S1(n8024));
    defparam sub_2032_add_2_33.INIT0 = 16'hf555;
    defparam sub_2032_add_2_33.INIT1 = 16'h0000;
    defparam sub_2032_add_2_33.INJECT1_0 = "NO";
    defparam sub_2032_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25621), .COUT(n25622));
    defparam sub_2032_add_2_31.INIT0 = 16'hf555;
    defparam sub_2032_add_2_31.INIT1 = 16'hf555;
    defparam sub_2032_add_2_31.INJECT1_0 = "NO";
    defparam sub_2032_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    CCU2D sub_2032_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25620), .COUT(n25621));
    defparam sub_2032_add_2_29.INIT0 = 16'hf555;
    defparam sub_2032_add_2_29.INIT1 = 16'hf555;
    defparam sub_2032_add_2_29.INJECT1_0 = "NO";
    defparam sub_2032_add_2_29.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n30300), .PD(n16223), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2032_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25619), .COUT(n25620));
    defparam sub_2032_add_2_27.INIT0 = 16'hf555;
    defparam sub_2032_add_2_27.INIT1 = 16'hf555;
    defparam sub_2032_add_2_27.INJECT1_0 = "NO";
    defparam sub_2032_add_2_27.INJECT1_1 = "NO";
    LUT4 i1021_2_lut_rep_291 (.A(n7990), .B(n32380), .Z(n30300)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1021_2_lut_rep_291.init = 16'heeee;
    FD1S3IX count_2614__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i1.GSR = "ENABLED";
    FD1S3IX count_2614__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i2.GSR = "ENABLED";
    FD1S3IX count_2614__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i3.GSR = "ENABLED";
    FD1S3IX count_2614__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i4.GSR = "ENABLED";
    FD1S3IX count_2614__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i5.GSR = "ENABLED";
    FD1S3IX count_2614__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i6.GSR = "ENABLED";
    FD1S3IX count_2614__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i7.GSR = "ENABLED";
    FD1S3IX count_2614__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i8.GSR = "ENABLED";
    FD1S3IX count_2614__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i9.GSR = "ENABLED";
    FD1S3IX count_2614__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i10.GSR = "ENABLED";
    FD1S3IX count_2614__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i11.GSR = "ENABLED";
    FD1S3IX count_2614__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i12.GSR = "ENABLED";
    FD1S3IX count_2614__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i13.GSR = "ENABLED";
    FD1S3IX count_2614__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i14.GSR = "ENABLED";
    FD1S3IX count_2614__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i15.GSR = "ENABLED";
    FD1S3IX count_2614__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i16.GSR = "ENABLED";
    FD1S3IX count_2614__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i17.GSR = "ENABLED";
    FD1S3IX count_2614__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i18.GSR = "ENABLED";
    FD1S3IX count_2614__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i19.GSR = "ENABLED";
    FD1S3IX count_2614__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i20.GSR = "ENABLED";
    FD1S3IX count_2614__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i21.GSR = "ENABLED";
    FD1S3IX count_2614__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i22.GSR = "ENABLED";
    FD1S3IX count_2614__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i23.GSR = "ENABLED";
    FD1S3IX count_2614__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i24.GSR = "ENABLED";
    FD1S3IX count_2614__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i25.GSR = "ENABLED";
    FD1S3IX count_2614__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i26.GSR = "ENABLED";
    FD1S3IX count_2614__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i27.GSR = "ENABLED";
    FD1S3IX count_2614__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i28.GSR = "ENABLED";
    FD1S3IX count_2614__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i29.GSR = "ENABLED";
    FD1S3IX count_2614__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i30.GSR = "ENABLED";
    FD1S3IX count_2614__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n30300), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614__i31.GSR = "ENABLED";
    CCU2D sub_2032_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25618), .COUT(n25619));
    defparam sub_2032_add_2_25.INIT0 = 16'hf555;
    defparam sub_2032_add_2_25.INIT1 = 16'hf555;
    defparam sub_2032_add_2_25.INJECT1_0 = "NO";
    defparam sub_2032_add_2_25.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n30300), .CD(n16223), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    LUT4 i9811_2_lut_3_lut (.A(n7990), .B(n32380), .C(n8024), .Z(n16223)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9811_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_2032_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25617), .COUT(n25618));
    defparam sub_2032_add_2_23.INIT0 = 16'hf555;
    defparam sub_2032_add_2_23.INIT1 = 16'hf555;
    defparam sub_2032_add_2_23.INJECT1_0 = "NO";
    defparam sub_2032_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25616), .COUT(n25617));
    defparam sub_2032_add_2_21.INIT0 = 16'hf555;
    defparam sub_2032_add_2_21.INIT1 = 16'hf555;
    defparam sub_2032_add_2_21.INJECT1_0 = "NO";
    defparam sub_2032_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25615), .COUT(n25616));
    defparam sub_2032_add_2_19.INIT0 = 16'hf555;
    defparam sub_2032_add_2_19.INIT1 = 16'hf555;
    defparam sub_2032_add_2_19.INJECT1_0 = "NO";
    defparam sub_2032_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25614), .COUT(n25615));
    defparam sub_2032_add_2_17.INIT0 = 16'hf555;
    defparam sub_2032_add_2_17.INIT1 = 16'hf555;
    defparam sub_2032_add_2_17.INJECT1_0 = "NO";
    defparam sub_2032_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25613), .COUT(n25614));
    defparam sub_2032_add_2_15.INIT0 = 16'hf555;
    defparam sub_2032_add_2_15.INIT1 = 16'hf555;
    defparam sub_2032_add_2_15.INJECT1_0 = "NO";
    defparam sub_2032_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25612), .COUT(n25613));
    defparam sub_2032_add_2_13.INIT0 = 16'hf555;
    defparam sub_2032_add_2_13.INIT1 = 16'hf555;
    defparam sub_2032_add_2_13.INJECT1_0 = "NO";
    defparam sub_2032_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26054), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_33.INIT1 = 16'h0000;
    defparam count_2614_add_4_33.INJECT1_0 = "NO";
    defparam count_2614_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26053), .COUT(n26054), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_31.INJECT1_0 = "NO";
    defparam count_2614_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25611), .COUT(n25612));
    defparam sub_2032_add_2_11.INIT0 = 16'hf555;
    defparam sub_2032_add_2_11.INIT1 = 16'hf555;
    defparam sub_2032_add_2_11.INJECT1_0 = "NO";
    defparam sub_2032_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26052), .COUT(n26053), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_29.INJECT1_0 = "NO";
    defparam count_2614_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26051), .COUT(n26052), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_27.INJECT1_0 = "NO";
    defparam count_2614_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25610), .COUT(n25611));
    defparam sub_2032_add_2_9.INIT0 = 16'hf555;
    defparam sub_2032_add_2_9.INIT1 = 16'hf555;
    defparam sub_2032_add_2_9.INJECT1_0 = "NO";
    defparam sub_2032_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25609), .COUT(n25610));
    defparam sub_2032_add_2_7.INIT0 = 16'hf555;
    defparam sub_2032_add_2_7.INIT1 = 16'hf555;
    defparam sub_2032_add_2_7.INJECT1_0 = "NO";
    defparam sub_2032_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2032_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25608), .COUT(n25609));
    defparam sub_2032_add_2_5.INIT0 = 16'hf555;
    defparam sub_2032_add_2_5.INIT1 = 16'hf555;
    defparam sub_2032_add_2_5.INJECT1_0 = "NO";
    defparam sub_2032_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26050), .COUT(n26051), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_25.INJECT1_0 = "NO";
    defparam count_2614_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26049), .COUT(n26050), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_23.INJECT1_0 = "NO";
    defparam count_2614_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2614_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26048), .COUT(n26049), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2614_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2614_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2614_add_4_21.INJECT1_0 = "NO";
    defparam count_2614_add_4_21.INJECT1_1 = "NO";
    
endmodule
