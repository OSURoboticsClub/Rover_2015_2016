// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Mon Apr 18 02:10:54 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(362[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    output expansion4 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[13:23])
    output expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(461[15:21])
    wire n33682 /* synthesis nomerge= */ ;
    
    wire GND_net, VCC_net, uart_rx_c, n10889, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, signal_light_c, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
        encoder_la_c, encoder_lb_c, encoder_li_c, rc_ch1_c, rc_ch2_c, 
        rc_ch3_c, rc_ch4_c, rc_ch7_c, rc_ch8_c, motor_pwm_l_c, xbee_pause_c, 
        debug_c_7, debug_c_5, debug_c_4, debug_c_3, debug_c_2, debug_c_0;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(457[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    
    wire rw, n14116, n27759, n27960, n14094;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(464[13:24])
    
    wire timeout_pause;
    wire [31:0]timeout_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[13:26])
    
    wire prev_uart_rx, clk_255kHz, n27887, n14258, n14374, n14372, 
        n1153, n31906, n5, n33685;
    wire [7:0]n8475;
    
    wire n154, n32;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n27769, n24, n27766, n8343, n34, n2954, n14369, n27768, 
        n8, n22, n27983;
    wire [31:0]n1468;
    
    wire n27877, n30466, n30426, n5811, n9198, n2863, n2853, n2850, 
        n13876;
    wire [31:0]n5951;
    
    wire n13557, n14358, n3984, n4, n5_adj_541, n30086, n3, n6, 
        n9362;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    
    wire clk_1Hz, prev_clk_1Hz;
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(32[12:21])
    
    wire prev_select, n46, n32_adj_542, n32_adj_543, n29174, n8_adj_544, 
        n6_adj_545, n4071;
    wire [7:0]\register[0]_adj_899 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [2:0]read_size_adj_901;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(93[12:21])
    
    wire n30445, n16566, n27226, n8_adj_547;
    wire [15:0]n281;
    
    wire n27225, n5_adj_548, n11158, n11020, n27224, n30220, n16565, 
        n241, n13797, n29175;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched, prev_limit_latched, step_clk, prev_step_clk;
    wire [31:0]read_value_adj_907;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_908;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_583, n27223, n27222, n27787, n8238, n27221, 
        n30196, n27220, n13779, n7, n8_adj_584, n21079, n13, n21082;
    wire [31:0]n580;
    
    wire n14, n22_adj_585, n13100, n2816;
    wire [7:0]control_reg_adj_916;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_917;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_918;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched_adj_587, prev_limit_latched_adj_588, int_step, 
        step_clk_adj_589, prev_step_clk_adj_590;
    wire [31:0]read_value_adj_919;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_920;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_625, n3_adj_626, n6_adj_627, n21084, n3_adj_628, 
        n3_adj_629, n6_adj_630, n8204, n13735, n22_adj_631, n6_adj_632, 
        n14661;
    wire [7:0]n5491;
    
    wire n110, n250, n13710, n13708, n13700, n13698, n111, n13693, 
        n29798, n29916;
    wire [7:0]control_reg_adj_957;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched_adj_634, prev_limit_latched_adj_635, step_clk_adj_636, 
        prev_step_clk_adj_637;
    wire [31:0]read_value_adj_960;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_961;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_672, n52, n3_adj_673, n3_adj_674, n6_adj_675, 
        n3_adj_676, n8134, n27886, n13667, n27883, n7892, n3_adj_677, 
        n31933, n9312, n9297;
    wire [31:0]n100_adj_1306;
    
    wire n29469, n12, n21092, n21090, n5_adj_679, n57, n46_adj_680, 
        n13647, n5_adj_681;
    wire [7:0]control_reg_adj_998;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched_adj_683, prev_limit_latched_adj_684;
    wire [31:0]read_value_adj_1001;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_1002;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_719, n13642, n29770, n8100;
    wire [31:0]n224_adj_1006;
    wire [31:0]n3899;
    
    wire n16545, n27853, n27809, n30202;
    wire [7:0]n571_adj_1020;
    
    wire n30166, n8_adj_724, n6_adj_725;
    wire [31:0]n99_adj_1308;
    wire [31:0]read_value_adj_1041;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[13:23])
    wire [2:0]read_size_adj_1042;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(67[12:21])
    
    wire prev_select_adj_760, n47, n13608, n3_adj_761, n6_adj_762;
    wire [31:0]read_value_adj_1048;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[13:23])
    wire [2:0]read_size_adj_1049;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(67[12:21])
    
    wire prev_select_adj_797, n1165, n14315, n6_adj_798, n3_adj_799, 
        n11927, n6_adj_800, n3_adj_801, n31928, n6_adj_802, n3_adj_803, 
        n6_adj_804, n3_adj_805, n6_adj_806;
    wire [14:0]n33921;
    
    wire n33687, n3_adj_814, n6_adj_815, n6_adj_816, n3_adj_817, n6_adj_818, 
        n94_adj_819, n6_adj_820, n31926, n33680, n31924, n31923, 
        n31922, n31921, n32090, n31920, n31919, n32089, n32088, 
        n31918, n3_adj_821, n6_adj_822, n11981, n33686, n31915, 
        n96_adj_823, n3_adj_824, n1, n27879, n3_adj_825, n6_adj_826, 
        n3_adj_827, n6_adj_828, n30361, n3_adj_829, n6_adj_830, n5_adj_831, 
        n8_adj_832, n4_adj_833, n8_adj_834, n42_adj_835, n5_adj_836, 
        n8_adj_837, n3_adj_838, n6_adj_839, n3_adj_840, n32080, n6_adj_841, 
        n40_adj_842, n22326;
    wire [3:0]n7645;
    wire [3:0]n33857;
    
    wire n38_adj_844, n8030, n36_adj_845, n34_adj_846, n22296, n30, 
        n29, n12_adj_847, n8_adj_848, n32075;
    wire [7:0]n8493;
    
    wire n26, n29900, n17, n16, n30381;
    wire [7:0]n8484;
    
    wire n15, n14519, n32074;
    wire [31:0]n6756;
    
    wire n26761, n30_adj_849, n31904, n16744, n29189;
    wire [3:0]state_adj_1082;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    
    wire select_clk, n32068;
    wire [31:0]n63_adj_1083;
    
    wire n31515, n27644, n32064, n6_adj_853, n9139, n32062, n8_adj_854, 
        n15_adj_855, n27956, n30378, n27757, n32056, n32053, n32052, 
        n26760, n27577, n28044, n3_adj_856, n29788, n29213;
    wire [1:0]n9_adj_1320;
    
    wire n25, n26_adj_858, n30_adj_859, n29_adj_860, n18379, n30510, 
        n32039, n1_adj_861, n7996, n4168, n32034, n7753;
    wire [31:0]n4401;
    
    wire n32032, n3_adj_862, n32030;
    wire [2:0]quadA_delayed_adj_1138;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [2:0]quadB_delayed_adj_1139;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n32025, n6_adj_863, n26759, n32016, n29198, n29212, n29214, 
        n29208, n29200, n29216, n29190, n29191, n29202, n31903, 
        n29210, n29204, n9366, n32011, n29192, n29194, n30505, 
        n29206, n32006, n29195, n29197, n29199, n29201, n26758, 
        n29203, n32005, n32004, n31911, n29205, n26757, n29207, 
        n29209, n29211, n29215, n32003, n29196, n29193, n30489, 
        n7718, n22230, n32001, n26756, n26755, n26754, n21480, 
        n26753;
    wire [15:0]count_adj_1167;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n26752, n26751, n5_adj_864, n27331, n27330, n22330, n31996, 
        n29948, n29341, n26750, n31991, n31990, n27329;
    wire [15:0]count_adj_1179;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n27328, n26749, n27327, n27326, n27325, n31987, n31986, 
        n29869, n31905, n29866, n27946, n29946, n27324, n27323, 
        n31982, n27322, n27321, n26748, n5_adj_867, n27, n18374, 
        n28, n29768, n31977, n30358, n31975, n5_adj_868, n5_adj_869, 
        n31972, n31970, n7926, n7683, n31910, n26747, n31965, 
        n31964, n47_adj_870, n31902, n31959, n33683, n31957, n31955, 
        n31953, n31952, n31951, n28101, n107, n31950;
    wire [3:0]state_adj_1228;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n27979, n31948, n30355, n31909, n31944, n13323, n31942, 
        n10962, n31940, n12930, n30512, n26746, n30514, n31938, 
        n1168, n31908, n30516, n30518, n1180, n31937, n31907, 
        n27758, n30520;
    
    VHI i2 (.Z(VCC_net));
    GlobalControlPeripheral global_control (.debug_c_c(debug_c_c), .n9312(n9312), 
            .n31991(n31991), .read_size({read_size}), .n14372(n14372), 
            .n27946(n27946), .\register[2][31] (\register[2] [31]), .\register[2][30] (\register[2] [30]), 
            .\register[2][29] (\register[2] [29]), .prev_clk_1Hz(prev_clk_1Hz), 
            .clk_1Hz(clk_1Hz), .\register[2][28] (\register[2] [28]), .\register[2][27] (\register[2] [27]), 
            .prev_select(prev_select), .\select[1] (select[1]), .\register[2][26] (\register[2] [26]), 
            .\register[2][25] (\register[2] [25]), .\register[2][24] (\register[2] [24]), 
            .\register[2][23] (\register[2] [23]), .\register[2][22] (\register[2] [22]), 
            .\register[2][21] (\register[2] [21]), .\register[2][20] (\register[2] [20]), 
            .\register[2][19] (\register[2] [19]), .\register[2][18] (\register[2] [18]), 
            .\register[2][17] (\register[2] [17]), .\register[2][16] (\register[2] [16]), 
            .\register[2][15] (\register[2] [15]), .\register[2][14] (\register[2] [14]), 
            .\register[2][13] (\register[2] [13]), .\register[2][12] (\register[2] [12]), 
            .\register[2][11] (\register[2] [11]), .\register[2][10] (\register[2] [10]), 
            .\register[2][9] (\register[2] [9]), .\register[2][8] (\register[2] [8]), 
            .\register[2][7] (\register[2] [7]), .\register[2][6] (\register[2] [6]), 
            .\register[2][5] (\register[2] [5]), .\register[2][4] (\register[2] [4]), 
            .\register[2][3] (\register[2] [3]), .rw(rw), .n46(n46), .n11158(n11158), 
            .\register_addr[1] (register_addr[1]), .\register_addr[0] (register_addr[0]), 
            .n32034(n32034), .\register_addr[5] (register_addr[5]), .n32032(n32032), 
            .\databus[1] (databus[1]), .timeout_pause(timeout_pause), .n32088(n32088), 
            .signal_light_c(signal_light_c), .\register[0][7] (\register[0]_adj_899 [7]), 
            .n32016(n32016), .n8(n8_adj_584), .n31937(n31937), .read_value({read_value}), 
            .n9362(n9362), .GND_net(GND_net), .xbee_pause_c(xbee_pause_c), 
            .n5980(n5951[3]), .n29197(n29197), .n29211(n29211), .n29213(n29213), 
            .n29207(n29207), .n29199(n29199), .n29215(n29215), .n29189(n29189), 
            .n29190(n29190), .n29201(n29201), .n29209(n29209), .n29203(n29203), 
            .n29191(n29191), .n29193(n29193), .n29205(n29205), .n29194(n29194), 
            .n29196(n29196), .n29198(n29198), .n29200(n29200), .n29202(n29202), 
            .n29204(n29204), .n29206(n29206), .n29208(n29208), .n29210(n29210), 
            .n250(n250), .n15(n15_adj_855), .n29214(n29214), .n29216(n29216), 
            .n29195(n29195), .n29192(n29192), .n31965(n31965), .n31975(n31975), 
            .n29212(n29212), .n32052(n32052), .n32005(n32005), .n31972(n31972), 
            .n2863(n2863), .n30358(n30358)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(520[45] 531[74])
    IFS1P3DX prev_uart_rx_58 (.D(uart_rx_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(prev_uart_rx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam prev_uart_rx_58.GSR = "ENABLED";
    FD1S3AX timeout_pause_60 (.D(n28101), .CK(debug_c_c), .Q(timeout_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_pause_60.GSR = "ENABLED";
    CCU2D add_30_15 (.A0(timeout_count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26752), .COUT(n26753), .S0(n100_adj_1306[13]), 
          .S1(n100_adj_1306[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_15.INIT0 = 16'h5aaa;
    defparam add_30_15.INIT1 = 16'h5aaa;
    defparam add_30_15.INJECT1_0 = "NO";
    defparam add_30_15.INJECT1_1 = "NO";
    VLO i1 (.Z(GND_net));
    CCU2D add_30_13 (.A0(timeout_count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26751), .COUT(n26752), .S0(n100_adj_1306[11]), 
          .S1(n100_adj_1306[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_13.INIT0 = 16'h5aaa;
    defparam add_30_13.INIT1 = 16'h5aaa;
    defparam add_30_13.INJECT1_0 = "NO";
    defparam add_30_13.INJECT1_1 = "NO";
    LUT4 i23200_4_lut (.A(n32064), .B(n5_adj_864), .C(n27983), .D(n27879), 
         .Z(n30512)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23200_4_lut.init = 16'h3233;
    FD1P3IX timeout_count__i0 (.D(n100_adj_1306[0]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i0.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n46_adj_680), .B(n30196), .C(n30202), .D(count_adj_1167[9]), 
         .Z(n29341)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i2_4_lut.init = 16'h0322;
    CCU2D add_30_11 (.A0(timeout_count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26750), .COUT(n26751), .S0(n100_adj_1306[9]), 
          .S1(n100_adj_1306[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_11.INIT0 = 16'h5aaa;
    defparam add_30_11.INIT1 = 16'h5aaa;
    defparam add_30_11.INJECT1_0 = "NO";
    defparam add_30_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(count_adj_1167[8]), .B(n32062), .C(count_adj_1167[5]), 
         .D(n27853), .Z(n46_adj_680)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'heaaa;
    LUT4 i22794_4_lut (.A(n27809), .B(n30086), .C(count_adj_1167[8]), 
         .D(n32080), .Z(n30202)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i22794_4_lut.init = 16'hfefc;
    LUT4 i8_2_lut (.A(timeout_count[1]), .B(timeout_count[4]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(timeout_count[6]), .B(n36_adj_845), .C(n26), .D(timeout_count[2]), 
         .Z(n40_adj_842)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i22682_2_lut (.A(count_adj_1167[6]), .B(count_adj_1167[7]), .Z(n30086)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22682_2_lut.init = 16'heeee;
    LUT4 i23202_4_lut_4_lut (.A(n1168), .B(n1180), .C(n29866), .D(n31964), 
         .Z(n30514)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+!(D))) */ ;
    defparam i23202_4_lut_4_lut.init = 16'hbb02;
    LUT4 i15693_4_lut (.A(n47_adj_870), .B(n13100), .C(n21480), .D(n29946), 
         .Z(n22296)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i15693_4_lut.init = 16'hfcec;
    LUT4 i23032_2_lut (.A(int_step), .B(control_reg_adj_916[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i23032_2_lut.init = 16'h9999;
    LUT4 i2_3_lut_rep_480 (.A(n22296), .B(reset_count[14]), .C(n7718), 
         .D(clk_255kHz), .Z(n33686)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_480.init = 16'h0080;
    LUT4 i2_3_lut (.A(reset_count[11]), .B(reset_count[12]), .C(reset_count[13]), 
         .Z(n13100)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(467[7:30])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i14886_2_lut (.A(reset_count[9]), .B(reset_count[10]), .Z(n21480)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14886_2_lut.init = 16'h8888;
    LUT4 Select_4247_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[7]), 
         .D(rw), .Z(n8_adj_834)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4247_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i15_2_lut_rep_342_3_lut (.A(select[3]), .B(n32030), .C(n33683), 
         .Z(n31959)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam i15_2_lut_rep_342_3_lut.init = 16'h8080;
    LUT4 Select_4192_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[26]), 
         .D(rw), .Z(n6_adj_818)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4192_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i114_2_lut_3_lut (.A(select[3]), .B(n32030), .C(prev_select_adj_797), 
         .Z(n14116)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam i114_2_lut_3_lut.init = 16'h0808;
    LUT4 Select_4248_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[6]), 
         .D(rw), .Z(n8_adj_832)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4248_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4249_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[5]), 
         .D(rw), .Z(n8_adj_837)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4249_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i29_2_lut_rep_436 (.A(uart_rx_c), .B(prev_uart_rx), .Z(n32053)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(481[7:29])
    defparam i29_2_lut_rep_436.init = 16'h6666;
    LUT4 Select_4250_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[4]), 
         .D(rw), .Z(n8_adj_854)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4250_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4251_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[3]), 
         .D(n33683), .Z(n8_adj_547)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4251_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4252_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[2]), 
         .D(n33683), .Z(n8)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4252_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4254_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[0]), 
         .D(n33683), .Z(n8_adj_724)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4254_i8_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4177_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[31]), 
         .D(n33683), .Z(n6_adj_806)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4177_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4180_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[30]), 
         .D(n33683), .Z(n6_adj_798)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4180_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4183_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[29]), 
         .D(n33683), .Z(n6_adj_800)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4183_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4186_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[28]), 
         .D(rw), .Z(n6_adj_545)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4186_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4189_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[27]), 
         .D(rw), .Z(n6_adj_822)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4189_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4195_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[25]), 
         .D(rw), .Z(n6_adj_816)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4195_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4216_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[18]), 
         .D(rw), .Z(n6_adj_675)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4216_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2711_2_lut_3_lut (.A(uart_rx_c), .B(prev_uart_rx), .C(n7683), 
         .Z(n9297)) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(481[7:29])
    defparam i2711_2_lut_3_lut.init = 16'h6f6f;
    CCU2D add_30_33 (.A0(timeout_count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26761), .S0(n100_adj_1306[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_33.INIT0 = 16'h5aaa;
    defparam add_30_33.INIT1 = 16'h0000;
    defparam add_30_33.INJECT1_0 = "NO";
    defparam add_30_33.INJECT1_1 = "NO";
    LUT4 Select_4213_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[19]), 
         .D(rw), .Z(n6_adj_762)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4213_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4210_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[20]), 
         .D(rw), .Z(n6_adj_632)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4210_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4207_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[21]), 
         .D(rw), .Z(n6_adj_820)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4207_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4204_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[22]), 
         .D(rw), .Z(n6_adj_804)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4204_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4201_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[23]), 
         .D(rw), .Z(n6_adj_802)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4201_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4198_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[24]), 
         .D(rw), .Z(n6_adj_815)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4198_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_rep_333_4_lut (.A(select[3]), .B(n32030), .C(n32011), 
         .D(prev_select_adj_797), .Z(n31950)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam i2_3_lut_rep_333_4_lut.init = 16'h0080;
    LUT4 i23155_4_lut (.A(n30466), .B(n17), .C(n15), .D(n16), .Z(n28101)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i23155_4_lut.init = 16'h8000;
    LUT4 Select_4219_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[17]), 
         .D(rw), .Z(n6_adj_630)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4219_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4222_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[16]), 
         .D(rw), .Z(n6_adj_863)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4222_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D add_30_31 (.A0(timeout_count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26760), .COUT(n26761), .S0(n100_adj_1306[29]), 
          .S1(n100_adj_1306[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_31.INIT0 = 16'h5aaa;
    defparam add_30_31.INIT1 = 16'h5aaa;
    defparam add_30_31.INJECT1_0 = "NO";
    defparam add_30_31.INJECT1_1 = "NO";
    LUT4 Select_4225_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[15]), 
         .D(rw), .Z(n6_adj_725)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4225_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4228_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[14]), 
         .D(rw), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4228_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4231_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[13]), 
         .D(rw), .Z(n6_adj_627)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4231_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4234_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[12]), 
         .D(rw), .Z(n6_adj_826)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4234_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4237_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[11]), 
         .D(rw), .Z(n6_adj_828)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4237_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4240_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[10]), 
         .D(rw), .Z(n6_adj_839)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4240_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4243_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[9]), 
         .D(rw), .Z(n6_adj_841)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4243_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4246_i6_2_lut_3_lut_4_lut (.A(select[3]), .B(n32030), .C(read_value_adj_1048[8]), 
         .D(rw), .Z(n6_adj_830)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4246_i6_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23110_2_lut_rep_374 (.A(n22296), .B(reset_count[14]), .Z(n31991)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i23110_2_lut_rep_374.init = 16'h7777;
    LUT4 i1_2_lut_rep_291_3_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), 
         .C(n8343), .D(select_clk), .Z(n31908)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_291_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1029_2_lut_rep_288_3_lut (.A(n22296), .B(reset_count[14]), .C(n7996), 
         .Z(n31905)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1029_2_lut_rep_288_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n8343), 
         .Z(n107)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i1033_2_lut_rep_285_3_lut (.A(n22296), .B(reset_count[14]), .C(n8100), 
         .Z(n31902)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1033_2_lut_rep_285_3_lut.init = 16'hf7f7;
    LUT4 i14693_2_lut_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n7718), 
         .Z(n241)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i14693_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i9914_2_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(n8030), 
         .D(n7996), .Z(n16545)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i9914_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i10142_2_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(n7926), 
         .D(n7892), .Z(n16744)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10142_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1_3_lut_4_lut_4_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), 
         .C(n31909), .D(state_adj_1082[0]), .Z(n33857[0])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i1_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h7f80;
    LUT4 i4_2_lut_rep_335_3_lut (.A(n22296), .B(reset_count[14]), .C(debug_c_0), 
         .Z(n31952)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i4_2_lut_rep_335_3_lut.init = 16'hf7f7;
    LUT4 i1_3_lut_rep_340_4_lut (.A(n22296), .B(reset_count[14]), .C(state_adj_1228[3]), 
         .D(state_adj_1228[2]), .Z(n31957)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_340_4_lut.init = 16'h0888;
    LUT4 i15028_2_lut_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(databus[0]), 
         .Z(n571_adj_1020[0])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15028_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_311_3_lut_4_lut (.A(n22296), .B(reset_count[14]), 
         .C(register_addr[1]), .D(register_addr[0]), .Z(n31928)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_311_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(prev_limit_latched_adj_684), 
         .D(limit_latched_adj_683), .Z(n11981)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h7f77;
    LUT4 i23184_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(state_adj_1228[2]), 
         .D(n31515), .Z(n14519)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i23184_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i4394_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(limit_latched_adj_634), 
         .D(prev_limit_latched_adj_635), .Z(n11020)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i4394_3_lut_4_lut.init = 16'h77f7;
    LUT4 i1_3_lut_4_lut_adj_474 (.A(n22296), .B(reset_count[14]), .C(prev_limit_latched), 
         .D(limit_latched), .Z(n10962)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_474.init = 16'h7f77;
    LUT4 i5301_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(limit_latched_adj_587), 
         .D(prev_limit_latched_adj_588), .Z(n11927)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i5301_3_lut_4_lut.init = 16'h77f7;
    LUT4 i23045_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n30355), 
         .Z(n2954)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i23045_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i23048_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n30358), 
         .Z(n2863)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i23048_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i23051_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n30361), 
         .Z(n2853)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i23051_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i972_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n7753), 
         .Z(n2816)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i972_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i23178_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n30489), 
         .Z(n22330)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i23178_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(n9139), .Z(n13698)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_adj_475 (.A(n22296), .B(reset_count[14]), .C(n13693), 
         .Z(n110)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_475.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_338_3_lut (.A(n22296), .B(reset_count[14]), .C(register_addr[0]), 
         .Z(n31955)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_338_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_476 (.A(n22296), .B(reset_count[14]), .C(n13667), 
         .Z(n111)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_476.init = 16'hf7f7;
    LUT4 i15417_2_lut_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(databus[7]), 
         .Z(n281[15])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15417_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_477 (.A(n22296), .B(reset_count[14]), .C(n13642), 
         .Z(n14258)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_477.init = 16'hf7f7;
    LUT4 i23075_2_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(n31926), 
         .D(register_addr[0]), .Z(n22326)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i23075_2_lut_3_lut_4_lut.init = 16'h77f7;
    CCU2D add_30_29 (.A0(timeout_count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26759), .COUT(n26760), .S0(n100_adj_1306[27]), 
          .S1(n100_adj_1306[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_29.INIT0 = 16'h5aaa;
    defparam add_30_29.INIT1 = 16'h5aaa;
    defparam add_30_29.INJECT1_0 = "NO";
    defparam add_30_29.INJECT1_1 = "NO";
    CCU2D add_30_27 (.A0(timeout_count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26758), .COUT(n26759), .S0(n100_adj_1306[25]), 
          .S1(n100_adj_1306[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_27.INIT0 = 16'h5aaa;
    defparam add_30_27.INIT1 = 16'h5aaa;
    defparam add_30_27.INJECT1_0 = "NO";
    defparam add_30_27.INJECT1_1 = "NO";
    LUT4 i9934_2_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(n8134), 
         .D(n8100), .Z(n16565)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i9934_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(n4401[0]), 
         .D(debug_c_0), .Z(n99_adj_1308[0])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i15481_2_lut_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(databus[4]), 
         .Z(n580[4])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15481_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i15477_2_lut_2_lut_3_lut (.A(n22296), .B(reset_count[14]), .C(databus[2]), 
         .Z(n580[2])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15477_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i2721_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(clk_1Hz), 
         .D(prev_clk_1Hz), .Z(n9312)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i2721_3_lut_4_lut.init = 16'h77f7;
    LUT4 i963_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(select[1]), 
         .D(prev_select), .Z(n14372)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i963_3_lut_4_lut.init = 16'h0080;
    LUT4 i2_3_lut_rep_289_4_lut (.A(n22296), .B(reset_count[14]), .C(n7718), 
         .D(clk_255kHz), .Z(n31906)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_289_4_lut.init = 16'h0080;
    LUT4 i1025_2_lut_rep_287_3_lut (.A(n22296), .B(reset_count[14]), .C(n7892), 
         .Z(n31904)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1025_2_lut_rep_287_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_4_lut_adj_478 (.A(n22296), .B(reset_count[14]), 
         .C(n31926), .D(register_addr[0]), .Z(n13557)) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_478.init = 16'hf777;
    LUT4 i9935_2_lut_3_lut_4_lut (.A(n22296), .B(reset_count[14]), .C(n8238), 
         .D(n8204), .Z(n16566)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i9935_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1037_2_lut_rep_286_3_lut (.A(n22296), .B(reset_count[14]), .C(n8204), 
         .Z(n31903)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1037_2_lut_rep_286_3_lut.init = 16'hf7f7;
    CCU2D reset_count_2631_2632_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27226), .S0(n33921[13]), 
          .S1(n33921[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2631_2632_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27225), .COUT(n27226), .S0(n33921[11]), 
          .S1(n33921[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2631_2632_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27224), .COUT(n27225), .S0(n33921[9]), 
          .S1(n33921[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2631_2632_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27223), .COUT(n27224), .S0(n33921[7]), 
          .S1(n33921[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2631_2632_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27222), .COUT(n27223), .S0(n33921[5]), 
          .S1(n33921[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_7.INJECT1_1 = "NO";
    CCU2D reset_count_2631_2632_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27221), .COUT(n27222), .S0(n33921[3]), 
          .S1(n33921[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_5.INJECT1_1 = "NO";
    CCU2D reset_count_2631_2632_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27220), .COUT(n27221), .S0(n33921[1]), 
          .S1(n33921[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2631_2632_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2631_2632_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27220), .S1(n33921[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2631_2632_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2631_2632_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2631_2632_add_4_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_479 (.A(n57), .B(n30220), .C(n154), .D(count_adj_1179[9]), 
         .Z(n29469)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i2_4_lut_adj_479.init = 16'h0322;
    LUT4 i1_2_lut (.A(count_adj_1179[8]), .B(n27644), .Z(n57)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i22812_4_lut (.A(count_adj_1179[13]), .B(count_adj_1179[10]), .C(count_adj_1179[11]), 
         .D(n32025), .Z(n30220)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22812_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_479 (.A(n22296), .B(reset_count[14]), .C(n7718), 
         .D(clk_255kHz), .Z(n33685)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_479.init = 16'h0080;
    LUT4 i23154_4_lut (.A(n29), .B(n42_adj_835), .C(n38_adj_844), .D(n30), 
         .Z(n30466)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i23154_4_lut.init = 16'h0001;
    LUT4 i23060_4_lut (.A(n29948), .B(reset_count[14]), .C(n13100), .D(n21480), 
         .Z(n30_adj_849)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i23060_4_lut.init = 16'h373f;
    LUT4 i1_4_lut_adj_480 (.A(n22230), .B(n29946), .C(reset_count[6]), 
         .D(reset_count[5]), .Z(n29948)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(471[17:42])
    defparam i1_4_lut_adj_480.init = 16'hfcec;
    LUT4 i15627_4_lut (.A(reset_count[0]), .B(reset_count[4]), .C(n6_adj_853), 
         .D(reset_count[3]), .Z(n22230)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i15627_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(reset_count[1]), .B(reset_count[2]), .Z(n6_adj_853)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_30_25 (.A0(timeout_count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26757), .COUT(n26758), .S0(n100_adj_1306[23]), 
          .S1(n100_adj_1306[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_25.INIT0 = 16'h5aaa;
    defparam add_30_25.INIT1 = 16'h5aaa;
    defparam add_30_25.INJECT1_0 = "NO";
    defparam add_30_25.INJECT1_1 = "NO";
    FD1P3AX reset_count_2631_2632__i1 (.D(n33921[0]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i1.GSR = "ENABLED";
    CCU2D add_30_23 (.A0(timeout_count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26756), .COUT(n26757), .S0(n100_adj_1306[21]), 
          .S1(n100_adj_1306[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_23.INIT0 = 16'h5aaa;
    defparam add_30_23.INIT1 = 16'h5aaa;
    defparam add_30_23.INJECT1_0 = "NO";
    defparam add_30_23.INJECT1_1 = "NO";
    LUT4 i15_2_lut_3_lut (.A(select[3]), .B(n32030), .C(rw), .Z(n47)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam i15_2_lut_3_lut.init = 16'h2020;
    LUT4 i114_2_lut_3_lut_adj_481 (.A(select[3]), .B(n32030), .C(prev_select_adj_760), 
         .Z(n13797)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam i114_2_lut_3_lut_adj_481.init = 16'h0202;
    LUT4 Select_4264_i8_2_lut_3_lut (.A(select[3]), .B(n32030), .C(read_size_adj_1042[0]), 
         .Z(n8_adj_544)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[4] 673[11])
    defparam Select_4264_i8_2_lut_3_lut.init = 16'h2020;
    CCU2D add_30_21 (.A0(timeout_count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26755), .COUT(n26756), .S0(n100_adj_1306[19]), 
          .S1(n100_adj_1306[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_21.INIT0 = 16'h5aaa;
    defparam add_30_21.INIT1 = 16'h5aaa;
    defparam add_30_21.INJECT1_0 = "NO";
    defparam add_30_21.INJECT1_1 = "NO";
    LUT4 i23198_4_lut (.A(n5_adj_867), .B(n32074), .C(n28044), .D(n27887), 
         .Z(n30510)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i23198_4_lut.init = 16'h5455;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n31991), .B(n29916), .C(n31933), .D(register_addr[0]), 
         .Z(n4168)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i2_3_lut_rep_481 (.A(n22296), .B(reset_count[14]), .C(n7718), 
         .D(clk_255kHz), .Z(n33687)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_481.init = 16'h0080;
    LUT4 i7_4_lut (.A(timeout_count[16]), .B(timeout_count[25]), .C(timeout_count[15]), 
         .D(timeout_count[24]), .Z(n17)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(timeout_count[8]), .B(timeout_count[20]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i6_4_lut (.A(timeout_count[17]), .B(timeout_count[9]), .C(timeout_count[23]), 
         .D(timeout_count[10]), .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i7_2_lut (.A(timeout_count[5]), .B(timeout_count[18]), .Z(n29)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(timeout_count[12]), .B(n40_adj_842), .C(n34_adj_846), 
         .D(timeout_count[19]), .Z(n42_adj_835)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_adj_482 (.A(reset_count[7]), .B(reset_count[5]), .C(reset_count[6]), 
         .Z(n27577)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_adj_482.init = 16'h8080;
    CCU2D add_30_9 (.A0(timeout_count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26749), .COUT(n26750), .S0(n100_adj_1306[7]), 
          .S1(n100_adj_1306[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_9.INIT0 = 16'h5aaa;
    defparam add_30_9.INIT1 = 16'h5aaa;
    defparam add_30_9.INJECT1_0 = "NO";
    defparam add_30_9.INJECT1_1 = "NO";
    LUT4 i16_4_lut (.A(timeout_count[31]), .B(timeout_count[22]), .C(timeout_count[21]), 
         .D(timeout_count[28]), .Z(n38_adj_844)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i16_4_lut.init = 16'hfffe;
    FD1P3IX timeout_count__i31 (.D(n100_adj_1306[31]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i31.GSR = "ENABLED";
    FD1P3IX timeout_count__i30 (.D(n100_adj_1306[30]), .SP(n9198), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i30.GSR = "ENABLED";
    FD1P3IX timeout_count__i29 (.D(n100_adj_1306[29]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i29.GSR = "ENABLED";
    FD1P3IX timeout_count__i28 (.D(n100_adj_1306[28]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i28.GSR = "ENABLED";
    FD1P3IX timeout_count__i27 (.D(n100_adj_1306[27]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i27.GSR = "ENABLED";
    FD1P3IX timeout_count__i26 (.D(n100_adj_1306[26]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i26.GSR = "ENABLED";
    FD1P3IX timeout_count__i25 (.D(n100_adj_1306[25]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i25.GSR = "ENABLED";
    FD1P3IX timeout_count__i24 (.D(n100_adj_1306[24]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i24.GSR = "ENABLED";
    FD1P3IX timeout_count__i23 (.D(n100_adj_1306[23]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i23.GSR = "ENABLED";
    FD1P3IX timeout_count__i22 (.D(n100_adj_1306[22]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i22.GSR = "ENABLED";
    FD1P3IX timeout_count__i21 (.D(n100_adj_1306[21]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i21.GSR = "ENABLED";
    FD1P3IX timeout_count__i20 (.D(n100_adj_1306[20]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i20.GSR = "ENABLED";
    FD1P3IX timeout_count__i19 (.D(n100_adj_1306[19]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i19.GSR = "ENABLED";
    FD1P3IX timeout_count__i18 (.D(n100_adj_1306[18]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i18.GSR = "ENABLED";
    FD1P3IX timeout_count__i17 (.D(n100_adj_1306[17]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i17.GSR = "ENABLED";
    FD1P3IX timeout_count__i16 (.D(n100_adj_1306[16]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i16.GSR = "ENABLED";
    FD1P3IX timeout_count__i15 (.D(n100_adj_1306[15]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i15.GSR = "ENABLED";
    FD1P3IX timeout_count__i14 (.D(n100_adj_1306[14]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i14.GSR = "ENABLED";
    FD1P3IX timeout_count__i13 (.D(n100_adj_1306[13]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i13.GSR = "ENABLED";
    FD1P3IX timeout_count__i12 (.D(n100_adj_1306[12]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i12.GSR = "ENABLED";
    FD1P3IX timeout_count__i11 (.D(n100_adj_1306[11]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i11.GSR = "ENABLED";
    FD1P3IX timeout_count__i10 (.D(n100_adj_1306[10]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i10.GSR = "ENABLED";
    FD1P3IX timeout_count__i9 (.D(n100_adj_1306[9]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i9.GSR = "ENABLED";
    FD1P3IX timeout_count__i8 (.D(n100_adj_1306[8]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i8.GSR = "ENABLED";
    FD1P3IX timeout_count__i7 (.D(n100_adj_1306[7]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i7.GSR = "ENABLED";
    FD1P3IX timeout_count__i6 (.D(n100_adj_1306[6]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i6.GSR = "ENABLED";
    FD1P3IX timeout_count__i5 (.D(n100_adj_1306[5]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i5.GSR = "ENABLED";
    FD1P3IX timeout_count__i4 (.D(n100_adj_1306[4]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i4.GSR = "ENABLED";
    FD1P3IX timeout_count__i3 (.D(n100_adj_1306[3]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i3.GSR = "ENABLED";
    FD1P3IX timeout_count__i2 (.D(n100_adj_1306[2]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i2.GSR = "ENABLED";
    FD1P3IX timeout_count__i1 (.D(n100_adj_1306[1]), .SP(n9297), .CD(n32053), 
            .CK(debug_c_c), .Q(timeout_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(478[9] 496[6])
    defparam timeout_count__i1.GSR = "ENABLED";
    CCU2D add_30_7 (.A0(timeout_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26748), .COUT(n26749), .S0(n100_adj_1306[5]), 
          .S1(n100_adj_1306[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_7.INIT0 = 16'h5aaa;
    defparam add_30_7.INIT1 = 16'h5aaa;
    defparam add_30_7.INJECT1_0 = "NO";
    defparam add_30_7.INJECT1_1 = "NO";
    LUT4 i12_4_lut (.A(timeout_count[14]), .B(timeout_count[11]), .C(timeout_count[30]), 
         .D(timeout_count[13]), .Z(n34_adj_846)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 Select_4253_i1_2_lut_3_lut_4_lut (.A(select[4]), .B(n31970), .C(read_value_adj_1001[1]), 
         .D(rw), .Z(n1_adj_861)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4253_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    PFUMX i11767 (.BLUT(n63_adj_1083[6]), .ALUT(n29_adj_860), .C0(n7), 
          .Z(n5491[6]));
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    IB encoder_li_pad (.I(encoder_li), .O(encoder_li_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    IB encoder_lb_pad (.I(encoder_lb), .O(encoder_lb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    IB encoder_la_pad (.I(encoder_la), .O(encoder_la_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    IB encoder_ri_pad (.I(encoder_ri), .O(encoder_ri_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    IB encoder_rb_pad (.I(encoder_rb), .O(encoder_rb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    IB encoder_ra_pad (.I(encoder_ra), .O(encoder_ra_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    LUT4 i1_2_lut_rep_294_3_lut_4_lut_4_lut (.A(select[4]), .B(n31970), 
         .C(n33683), .D(prev_select_adj_719), .Z(n31911)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_294_3_lut_4_lut_4_lut.init = 16'h0008;
    IB uart_rx_pad (.I(uart_rx), .O(uart_rx_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    OB debug_pad_0 (.I(debug_c_0), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_1 (.I(n10889), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_6 (.I(n31991), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB motor_pwm_r_pad (.I(GND_net), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    OB expansion5_pad (.I(GND_net), .O(expansion5));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    OB expansion4_pad (.I(GND_net), .O(expansion4));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[13:23])
    OB expansion3_pad (.I(GND_net), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion2_pad (.I(GND_net), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB expansion1_pad (.I(GND_net), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    LUT4 i14_4_lut (.A(timeout_count[29]), .B(timeout_count[26]), .C(timeout_count[7]), 
         .D(timeout_count[3]), .Z(n36_adj_845)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i14_4_lut.init = 16'hfffe;
    PFUMX i11747 (.BLUT(n63_adj_1083[3]), .ALUT(n25), .C0(n7), .Z(n18374));
    LUT4 i1_2_lut_adj_483 (.A(register_addr[4]), .B(register_addr[5]), .Z(n13323)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(552[4] 581[11])
    defparam i1_2_lut_adj_483.init = 16'h8888;
    PFUMX i11752 (.BLUT(n63_adj_1083[1]), .ALUT(n27), .C0(n7), .Z(n18379));
    PFUMX i11757 (.BLUT(n63_adj_1083[2]), .ALUT(n26_adj_858), .C0(n7), 
          .Z(n5491[2]));
    LUT4 i4_2_lut (.A(timeout_count[0]), .B(timeout_count[27]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(491[7:35])
    defparam i4_2_lut.init = 16'heeee;
    PFUMX i11762 (.BLUT(n63_adj_1083[4]), .ALUT(n28), .C0(n7), .Z(n5491[4]));
    PFUMX i11772 (.BLUT(n63_adj_1083[5]), .ALUT(n30_adj_859), .C0(n7), 
          .Z(n5491[5]));
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB uart_tx_pad (.I(n10889), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    CCU2D add_30_19 (.A0(timeout_count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26754), .COUT(n26755), .S0(n100_adj_1306[17]), 
          .S1(n100_adj_1306[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_19.INIT0 = 16'h5aaa;
    defparam add_30_19.INIT1 = 16'h5aaa;
    defparam add_30_19.INJECT1_0 = "NO";
    defparam add_30_19.INJECT1_1 = "NO";
    FD1P3AX reset_count_2631_2632__i2 (.D(n33921[1]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i2.GSR = "ENABLED";
    LUT4 i2621_1_lut (.A(n7683), .Z(n9198)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2621_1_lut.init = 16'h5555;
    LUT4 i14494_3_lut (.A(Stepper_Y_Dir_c), .B(div_factor_reg_adj_917[5]), 
         .C(register_addr[1]), .Z(n21090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    defparam i14494_3_lut.init = 16'hcaca;
    CCU2D add_30_17 (.A0(timeout_count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26753), .COUT(n26754), .S0(n100_adj_1306[15]), 
          .S1(n100_adj_1306[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_17.INIT0 = 16'h5aaa;
    defparam add_30_17.INIT1 = 16'h5aaa;
    defparam add_30_17.INJECT1_0 = "NO";
    defparam add_30_17.INJECT1_1 = "NO";
    LUT4 i14486_3_lut (.A(Stepper_Y_En_c), .B(div_factor_reg_adj_917[6]), 
         .C(register_addr[1]), .Z(n21082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    defparam i14486_3_lut.init = 16'hcaca;
    LUT4 i14483_3_lut (.A(control_reg_adj_916[3]), .B(div_factor_reg_adj_917[3]), 
         .C(register_addr[1]), .Z(n21079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    defparam i14483_3_lut.init = 16'hcaca;
    CCU2D add_30_5 (.A0(timeout_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26747), .COUT(n26748), .S0(n100_adj_1306[3]), 
          .S1(n100_adj_1306[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_5.INIT0 = 16'h5aaa;
    defparam add_30_5.INIT1 = 16'h5aaa;
    defparam add_30_5.INJECT1_0 = "NO";
    defparam add_30_5.INJECT1_1 = "NO";
    CCU2D add_30_3 (.A0(timeout_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26746), .COUT(n26747), .S0(n100_adj_1306[1]), 
          .S1(n100_adj_1306[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_3.INIT0 = 16'h5aaa;
    defparam add_30_3.INIT1 = 16'h5aaa;
    defparam add_30_3.INJECT1_0 = "NO";
    defparam add_30_3.INJECT1_1 = "NO";
    CCU2D add_30_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(timeout_count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26746), .S1(n100_adj_1306[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(488[24:41])
    defparam add_30_1.INIT0 = 16'hF000;
    defparam add_30_1.INIT1 = 16'h5555;
    defparam add_30_1.INJECT1_0 = "NO";
    defparam add_30_1.INJECT1_1 = "NO";
    FD1P3AX reset_count_2631_2632__i3 (.D(n33921[2]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i4 (.D(n33921[3]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i5 (.D(n33921[4]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i6 (.D(n33921[5]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i7 (.D(n33921[6]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i8 (.D(n33921[7]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i9 (.D(n33921[8]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i10 (.D(n33921[9]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i11 (.D(n33921[10]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i12 (.D(n33921[11]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i13 (.D(n33921[12]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i14 (.D(n33921[13]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2631_2632__i15 (.D(n33921[14]), .SP(n30_adj_849), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[20:35])
    defparam reset_count_2631_2632__i15.GSR = "ENABLED";
    PFUMX i14496 (.BLUT(n21090), .ALUT(n14), .C0(register_addr[0]), .Z(n21092));
    PFUMX i14488 (.BLUT(n21082), .ALUT(n13), .C0(register_addr[0]), .Z(n21084));
    PFUMX i14485 (.BLUT(n21079), .ALUT(n12), .C0(register_addr[0]), .Z(n6756[3]));
    CCU2D add_20098_24 (.A0(timeout_count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27331), .S1(n7683));
    defparam add_20098_24.INIT0 = 16'h5555;
    defparam add_20098_24.INIT1 = 16'h0000;
    defparam add_20098_24.INJECT1_0 = "NO";
    defparam add_20098_24.INJECT1_1 = "NO";
    CCU2D add_20098_22 (.A0(timeout_count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27330), .COUT(n27331));
    defparam add_20098_22.INIT0 = 16'h5555;
    defparam add_20098_22.INIT1 = 16'h5555;
    defparam add_20098_22.INJECT1_0 = "NO";
    defparam add_20098_22.INJECT1_1 = "NO";
    CCU2D add_20098_20 (.A0(timeout_count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27329), .COUT(n27330));
    defparam add_20098_20.INIT0 = 16'h5555;
    defparam add_20098_20.INIT1 = 16'h5555;
    defparam add_20098_20.INJECT1_0 = "NO";
    defparam add_20098_20.INJECT1_1 = "NO";
    CCU2D add_20098_18 (.A0(timeout_count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27328), .COUT(n27329));
    defparam add_20098_18.INIT0 = 16'h5aaa;
    defparam add_20098_18.INIT1 = 16'h5555;
    defparam add_20098_18.INJECT1_0 = "NO";
    defparam add_20098_18.INJECT1_1 = "NO";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2D add_20098_16 (.A0(timeout_count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27327), .COUT(n27328));
    defparam add_20098_16.INIT0 = 16'h5aaa;
    defparam add_20098_16.INIT1 = 16'h5aaa;
    defparam add_20098_16.INJECT1_0 = "NO";
    defparam add_20098_16.INJECT1_1 = "NO";
    CCU2D add_20098_14 (.A0(timeout_count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27326), .COUT(n27327));
    defparam add_20098_14.INIT0 = 16'h5555;
    defparam add_20098_14.INIT1 = 16'h5555;
    defparam add_20098_14.INJECT1_0 = "NO";
    defparam add_20098_14.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_484 (.A(div_factor_reg_adj_917[9]), .B(n29770), .C(steps_reg_adj_918[9]), 
         .D(register_addr[0]), .Z(n29788)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    defparam i1_4_lut_adj_484.init = 16'hc088;
    CCU2D add_20098_12 (.A0(timeout_count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27325), .COUT(n27326));
    defparam add_20098_12.INIT0 = 16'h5555;
    defparam add_20098_12.INIT1 = 16'h5aaa;
    defparam add_20098_12.INJECT1_0 = "NO";
    defparam add_20098_12.INJECT1_1 = "NO";
    EncoderPeripheral_U11 left_encoder (.\read_size[0] (read_size_adj_1042[0]), 
            .debug_c_c(debug_c_c), .n13797(n13797), .n31923(n31923), .n27946(n27946), 
            .prev_select(prev_select_adj_760), .n32001(n32001), .read_value({read_value_adj_1041}), 
            .\read_size[2] (read_size_adj_1042[2]), .n15(n15_adj_855), .\register_addr[0] (register_addr[0]), 
            .n31952(n31952), .\quadA_delayed[2] (quadA_delayed_adj_1138[2]), 
            .\quadB_delayed[1] (quadB_delayed_adj_1139[1]), .n13779(n13779), 
            .encoder_li_c(encoder_li_c), .encoder_lb_c(encoder_lb_c), .encoder_la_c(encoder_la_c), 
            .VCC_net(VCC_net), .GND_net(GND_net), .\quadA_delayed[1] (quadA_delayed_adj_1138[1]), 
            .\quadB_delayed[2] (quadB_delayed_adj_1139[2])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(675[20] 685[47])
    CCU2D add_20098_10 (.A0(timeout_count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27324), .COUT(n27325));
    defparam add_20098_10.INIT0 = 16'h5aaa;
    defparam add_20098_10.INIT1 = 16'h5555;
    defparam add_20098_10.INJECT1_0 = "NO";
    defparam add_20098_10.INJECT1_1 = "NO";
    CCU2D add_20098_8 (.A0(timeout_count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27323), .COUT(n27324));
    defparam add_20098_8.INIT0 = 16'h5aaa;
    defparam add_20098_8.INIT1 = 16'h5aaa;
    defparam add_20098_8.INJECT1_0 = "NO";
    defparam add_20098_8.INJECT1_1 = "NO";
    CCU2D add_20098_6 (.A0(timeout_count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27322), .COUT(n27323));
    defparam add_20098_6.INIT0 = 16'h5555;
    defparam add_20098_6.INIT1 = 16'h5555;
    defparam add_20098_6.INJECT1_0 = "NO";
    defparam add_20098_6.INJECT1_1 = "NO";
    CCU2D add_20098_4 (.A0(timeout_count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27321), .COUT(n27322));
    defparam add_20098_4.INIT0 = 16'h5555;
    defparam add_20098_4.INIT1 = 16'h5555;
    defparam add_20098_4.INJECT1_0 = "NO";
    defparam add_20098_4.INJECT1_1 = "NO";
    CCU2D add_20098_2 (.A0(timeout_count[9]), .B0(timeout_count[8]), .C0(GND_net), 
          .D0(GND_net), .A1(timeout_count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27321));
    defparam add_20098_2.INIT0 = 16'h7000;
    defparam add_20098_2.INIT1 = 16'h5aaa;
    defparam add_20098_2.INJECT1_0 = "NO";
    defparam add_20098_2.INJECT1_1 = "NO";
    RCPeripheral rc_receiver (.databus_out({databus_out}), .n33683(n33683), 
            .read_value({read_value_adj_960}), .read_value_adj_264({read_value}), 
            .n52(n52), .n46(n46), .n3(n3_adj_628), .databus({databus}), 
            .\read_value[16]_adj_83 (read_value_adj_1001[16]), .read_value_adj_265({read_value_adj_1041}), 
            .n31924(n31924), .n47(n47), .\read_value[16]_adj_116 (read_value_adj_907[16]), 
            .n6(n6_adj_863), .n31942(n31942), .n3_adj_117(n3_adj_856), 
            .\read_value[15]_adj_118 (read_value_adj_1001[15]), .\read_value[15]_adj_119 (read_value_adj_907[15]), 
            .n6_adj_120(n6_adj_725), .rw(rw), .\register_addr[0] (register_addr[0]), 
            .n3_adj_121(n3), .\read_value[14]_adj_122 (read_value_adj_1001[14]), 
            .\read_value[14]_adj_123 (read_value_adj_907[14]), .n6_adj_124(n6), 
            .\select[7] (select[7]), .n3_adj_125(n3_adj_862), .\read_value[13]_adj_126 (read_value_adj_1001[13]), 
            .\read_value[13]_adj_127 (read_value_adj_907[13]), .n6_adj_128(n6_adj_627), 
            .n3_adj_129(n3_adj_799), .\read_value[30]_adj_130 (read_value_adj_1001[30]), 
            .\read_value[30]_adj_131 (read_value_adj_907[30]), .n6_adj_132(n6_adj_798), 
            .n3_adj_133(n3_adj_825), .\read_value[12]_adj_134 (read_value_adj_1001[12]), 
            .\read_value[12]_adj_135 (read_value_adj_907[12]), .n6_adj_136(n6_adj_826), 
            .n3_adj_137(n3_adj_801), .\read_value[29]_adj_138 (read_value_adj_1001[29]), 
            .\read_value[29]_adj_139 (read_value_adj_907[29]), .n6_adj_140(n6_adj_800), 
            .n3_adj_141(n3_adj_626), .\read_value[28]_adj_142 (read_value_adj_1001[28]), 
            .\read_value[28]_adj_143 (read_value_adj_907[28]), .n6_adj_144(n6_adj_545), 
            .n3_adj_145(n3_adj_821), .\read_value[27]_adj_146 (read_value_adj_1001[27]), 
            .\read_value[27]_adj_147 (read_value_adj_907[27]), .n6_adj_148(n6_adj_822), 
            .n3_adj_149(n3_adj_827), .\read_value[11]_adj_150 (read_value_adj_1001[11]), 
            .\read_value[11]_adj_151 (read_value_adj_907[11]), .n6_adj_152(n6_adj_828), 
            .\register_addr[2] (register_addr[2]), .n3_adj_153(n3_adj_817), 
            .\read_value[26]_adj_154 (read_value_adj_1001[26]), .\read_value[26]_adj_155 (read_value_adj_907[26]), 
            .n6_adj_156(n6_adj_818), .n3_adj_157(n3_adj_838), .\read_value[10]_adj_158 (read_value_adj_1001[10]), 
            .\read_value[10]_adj_159 (read_value_adj_907[10]), .n6_adj_160(n6_adj_839), 
            .\read_value[0]_adj_161 (read_value_adj_919[0]), .n31944(n31944), 
            .n3_adj_162(n3_adj_840), .\read_value[9]_adj_163 (read_value_adj_1001[9]), 
            .\read_value[9]_adj_164 (read_value_adj_907[9]), .n6_adj_165(n6_adj_841), 
            .\read_value[0]_adj_166 (read_value_adj_907[0]), .read_size({read_size}), 
            .\select[1] (select[1]), .n32068(n32068), .\sendcount[1] (sendcount[1]), 
            .n12930(n12930), .n3_adj_167(n3_adj_829), .\read_value[8]_adj_168 (read_value_adj_1001[8]), 
            .n3_adj_169(n3_adj_677), .\read_value[25]_adj_170 (read_value_adj_1001[25]), 
            .\read_value[25]_adj_171 (read_value_adj_907[25]), .n6_adj_172(n6_adj_816), 
            .\read_value[8]_adj_173 (read_value_adj_907[8]), .n6_adj_174(n6_adj_830), 
            .\read_value[7]_adj_175 (read_value_adj_1001[7]), .n5(n5_adj_541), 
            .n8(n8_adj_834), .n3_adj_176(n3_adj_814), .\read_value[24]_adj_177 (read_value_adj_1001[24]), 
            .\read_value[24]_adj_178 (read_value_adj_907[24]), .n6_adj_179(n6_adj_815), 
            .\register_addr[1] (register_addr[1]), .\read_value[7]_adj_180 (read_value_adj_919[7]), 
            .\read_value[7]_adj_181 (read_value_adj_907[7]), .n3_adj_182(n3_adj_803), 
            .\read_value[23]_adj_183 (read_value_adj_1001[23]), .\read_value[23]_adj_184 (read_value_adj_907[23]), 
            .n6_adj_185(n6_adj_802), .n3_adj_186(n3_adj_676), .\read_value[22]_adj_187 (read_value_adj_1001[22]), 
            .\read_value[22]_adj_188 (read_value_adj_907[22]), .n6_adj_189(n6_adj_804), 
            .n3_adj_190(n3_adj_824), .\read_value[21]_adj_191 (read_value_adj_1001[21]), 
            .\read_value[21]_adj_192 (read_value_adj_907[21]), .n6_adj_193(n6_adj_820), 
            .n3_adj_194(n3_adj_673), .\read_value[20]_adj_195 (read_value_adj_1001[20]), 
            .\read_value[20]_adj_196 (read_value_adj_907[20]), .n6_adj_197(n6_adj_632), 
            .n3_adj_198(n3_adj_761), .\read_value[19]_adj_199 (read_value_adj_1001[19]), 
            .\read_value[19]_adj_200 (read_value_adj_907[19]), .n6_adj_201(n6_adj_762), 
            .n32090(n32090), .\register_addr[3] (register_addr[3]), .n32089(n32089), 
            .n31987(n31987), .n13323(n13323), .n31970(n31970), .\register_addr[5] (register_addr[5]), 
            .n31972(n31972), .n33680(n33680), .n31975(n31975), .n3_adj_202(n3_adj_674), 
            .n32034(n32034), .n32006(n32006), .\read_value[18]_adj_203 (read_value_adj_1001[18]), 
            .\read_value[18]_adj_204 (read_value_adj_907[18]), .n6_adj_205(n6_adj_675), 
            .n31965(n31965), .\select[4] (select[4]), .\read_size[0]_adj_206 (read_size_adj_1002[0]), 
            .n22(n22_adj_631), .\read_size[0]_adj_207 (read_size_adj_901[0]), 
            .n8_adj_208(n8_adj_544), .\select[2] (select[2]), .n12(n12_adj_847), 
            .n31990(n31990), .\read_size[0]_adj_209 (read_size_adj_1049[0]), 
            .n8_adj_210(n8_adj_848), .\read_size[0]_adj_211 (read_size_adj_908[0]), 
            .n30166(n30166), .\read_size[0]_adj_212 (read_size_adj_961[0]), 
            .n31977(n31977), .\read_size[0]_adj_213 (read_size_adj_920[0]), 
            .n3_adj_214(n3_adj_629), .\read_value[17]_adj_215 (read_value_adj_1001[17]), 
            .\read_value[17]_adj_216 (read_value_adj_907[17]), .n6_adj_217(n6_adj_630), 
            .\reg_size[2] (reg_size[2]), .\read_size[2]_adj_218 (read_size_adj_1042[2]), 
            .n32001(n32001), .\read_size[2]_adj_219 (read_size_adj_920[2]), 
            .\read_size[2]_adj_220 (read_size_adj_1049[2]), .\read_size[2]_adj_221 (read_size_adj_1002[2]), 
            .\read_size[2]_adj_222 (read_size_adj_908[2]), .\read_size[2]_adj_223 (read_size_adj_961[2]), 
            .\read_value[6]_adj_224 (read_value_adj_1001[6]), .n5_adj_225(n5_adj_831), 
            .n8_adj_226(n8_adj_832), .\read_value[6]_adj_227 (read_value_adj_919[6]), 
            .n4(n4), .\read_value[6]_adj_228 (read_value_adj_907[6]), .\read_value[1]_adj_229 (read_value_adj_1048[1]), 
            .n31959(n31959), .\read_value[5]_adj_230 (read_value_adj_1001[5]), 
            .n5_adj_231(n5_adj_836), .n8_adj_232(n8_adj_837), .\read_value[5]_adj_233 (read_value_adj_919[5]), 
            .\read_value[5]_adj_234 (read_value_adj_907[5]), .n32004(n32004), 
            .\read_value[4]_adj_235 (read_value_adj_1001[4]), .n5_adj_236(n5_adj_869), 
            .n1(n1_adj_861), .n5_adj_237(n5_adj_679), .n8_adj_238(n8_adj_854), 
            .\read_value[4]_adj_239 (read_value_adj_919[4]), .\read_value[4]_adj_240 (read_value_adj_907[4]), 
            .\read_value[3]_adj_241 (read_value_adj_1001[3]), .n5_adj_242(n5), 
            .n8_adj_243(n8_adj_547), .\read_value[3]_adj_244 (read_value_adj_919[3]), 
            .\read_value[3]_adj_245 (read_value_adj_907[3]), .\read_value[2]_adj_246 (read_value_adj_1001[2]), 
            .n5_adj_247(n5_adj_548), .\read_value[1]_adj_248 (read_value_adj_919[1]), 
            .n3_adj_249(n3_adj_805), .\read_value[31]_adj_250 (read_value_adj_1001[31]), 
            .\read_value[31]_adj_251 (read_value_adj_907[31]), .n6_adj_252(n6_adj_806), 
            .n8_adj_253(n8), .\read_value[2]_adj_254 (read_value_adj_919[2]), 
            .\read_value[0]_adj_255 (read_value_adj_1001[0]), .n5_adj_256(n5_adj_681), 
            .\read_value[2]_adj_257 (read_value_adj_907[2]), .n8_adj_258(n8_adj_724), 
            .n32039(n32039), .n5_adj_259(n5_adj_868), .n27979(n27979), 
            .GND_net(GND_net), .debug_c_c(debug_c_c), .n33686(n33686), 
            .rc_ch8_c(rc_ch8_c), .n30381(n30381), .n33685(n33685), .n13735(n13735), 
            .n27956(n27956), .n27877(n27877), .rc_ch7_c(rc_ch7_c), .n5_adj_260(n5_adj_867), 
            .n32074(n32074), .n28044(n28044), .n27887(n27887), .n27759(n27759), 
            .n33687(n33687), .n14315(n14315), .n30505(n30505), .\count[8] (count_adj_1179[8]), 
            .\count[13] (count_adj_1179[13]), .n27644(n27644), .rc_ch4_c(rc_ch4_c), 
            .\count[11] (count_adj_1179[11]), .n30520(n30520), .\count[9] (count_adj_1179[9]), 
            .\count[10] (count_adj_1179[10]), .n32025(n32025), .n154(n154), 
            .n27883(n27883), .n29469(n29469), .n30220(n30220), .n5_adj_261(n5_adj_864), 
            .n27879(n27879), .n30196(n30196), .n27809(n27809), .\count[8]_adj_262 (count_adj_1167[8]), 
            .n30202(n30202), .\count[9]_adj_263 (count_adj_1167[9]), .\count[6] (count_adj_1167[6]), 
            .\count[7] (count_adj_1167[7]), .n32062(n32062), .\count[5] (count_adj_1167[5]), 
            .n27853(n27853), .n32064(n32064), .n27983(n27983), .rc_ch3_c(rc_ch3_c), 
            .n32080(n32080), .n27758(n27758), .n29341(n29341), .n14358(n14358), 
            .n30445(n30445), .n1168(n1168), .n1180(n1180), .n31964(n31964), 
            .n30426(n30426), .n31906(n31906), .n14369(n14369), .n27757(n27757), 
            .rc_ch2_c(rc_ch2_c), .n29866(n29866), .n1153(n1153), .n1165(n1165), 
            .n31948(n31948), .n30378(n30378), .n14374(n14374), .rc_ch1_c(rc_ch1_c), 
            .n27960(n27960), .n29869(n29869)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(699[15] 711[41])
    SabertoothSerialPeripheral motor_serial (.debug_c_c(debug_c_c), .n13557(n13557), 
            .n282(n281[15]), .n31991(n31991), .\databus[6] (databus[6]), 
            .\databus[5] (databus[5]), .\databus[4] (databus[4]), .\databus[3] (databus[3]), 
            .\databus[2] (databus[2]), .\databus[1] (databus[1]), .\databus[0] (databus[0]), 
            .\register[0] ({\register[0]_adj_899 [7], Open_0, Open_1, 
            Open_2, Open_3, Open_4, Open_5, Open_6}), .n22326(n22326), 
            .\read_size[0] (read_size_adj_901[0]), .n31922(n31922), .\select[2] (select[2]), 
            .n9366(n9366), .rw(rw), .n32075(n32075), .n31940(n31940), 
            .\register_addr[0] (register_addr[0]), .\reset_count[14] (reset_count[14]), 
            .n22296(n22296), .n5(n5_adj_541), .n5_adj_44(n5_adj_831), 
            .n5_adj_45(n5_adj_836), .n5_adj_46(n5_adj_869), .n5_adj_47(n5), 
            .n5_adj_48(n5_adj_681), .n5_adj_49(n5_adj_679), .n32088(n32088), 
            .n89(n63_adj_1083[6]), .n5_adj_50(n5_adj_548), .\state[0] (state_adj_1082[0]), 
            .GND_net(GND_net), .n12(n33857[0]), .n31907(n31907), .n7(n7), 
            .n31908(n31908), .n18379(n18379), .n5497(n5491[2]), .n18374(n18374), 
            .n5495(n5491[4]), .n5494(n5491[5]), .n5493(n5491[6]), .n32016(n32016), 
            .n29(n29_adj_860), .\state[1] (state_adj_1082[1]), .n7648(n7645[1]), 
            .n92(n63_adj_1083[3]), .n25(n25), .n94(n63_adj_1083[1]), .n27(n27), 
            .n93(n63_adj_1083[2]), .n26(n26_adj_858), .n91(n63_adj_1083[4]), 
            .n28(n28), .n90(n63_adj_1083[5]), .n30(n30_adj_859), .\reset_count[6] (reset_count[6]), 
            .\reset_count[5] (reset_count[5]), .\reset_count[4] (reset_count[4]), 
            .n47(n47_adj_870), .\reset_count[8] (reset_count[8]), .\reset_count[7] (reset_count[7]), 
            .n29946(n29946), .\state[3] (state_adj_1228[3]), .\state[2] (state_adj_1228[2]), 
            .n31515(n31515), .\reset_count[11] (reset_count[11]), .n21480(n21480), 
            .n27577(n27577), .n29900(n29900), .n14519(n14519), .n31957(n31957), 
            .motor_pwm_l_c(motor_pwm_l_c), .n8343(n8343), .n2954(n2954), 
            .n30355(n30355), .select_clk(select_clk), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(534[29] 542[56])
    LUT4 i2_3_lut_4_lut_4_lut_adj_485 (.A(n31991), .B(n32075), .C(n31975), 
         .D(register_addr[1]), .Z(n9366)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut_adj_485.init = 16'h4440;
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 i2_3_lut_3_lut (.A(n31996), .B(n1468[17]), .C(n1468[20]), .Z(n27886)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i2_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i23072_4_lut_4_lut (.A(n31996), .B(n4_adj_833), .C(n5811), .D(n1468[14]), 
         .Z(n13608)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i23072_4_lut_4_lut.init = 16'h2a00;
    LUT4 i23206_4_lut (.A(n32039), .B(n5_adj_868), .C(n27979), .D(n27877), 
         .Z(n30518)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23206_4_lut.init = 16'h3233;
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.debug_c_c(debug_c_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .n31991(n31991), .\read_size[0] (read_size_adj_920[0]), .n13700(n13700), 
            .n96(n96_adj_823), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), .n111(n111), 
            .n579(n571_adj_1020[0]), .prev_step_clk(prev_step_clk_adj_590), 
            .step_clk(step_clk_adj_589), .limit_latched(limit_latched_adj_587), 
            .prev_limit_latched(prev_limit_latched_adj_588), .n14094(n14094), 
            .prev_select(prev_select_adj_625), .n31977(n31977), .\register_addr[0] (register_addr[0]), 
            .\register_addr[1] (register_addr[1]), .n27769(n27769), .n31953(n31953), 
            .databus({databus}), .\div_factor_reg[9] (div_factor_reg_adj_917[9]), 
            .\div_factor_reg[6] (div_factor_reg_adj_917[6]), .\div_factor_reg[5] (div_factor_reg_adj_917[5]), 
            .\div_factor_reg[3] (div_factor_reg_adj_917[3]), .\control_reg[7] (control_reg_adj_916[7]), 
            .n13667(n13667), .n11927(n11927), .Stepper_Y_En_c(Stepper_Y_En_c), 
            .Stepper_Y_Dir_c(Stepper_Y_Dir_c), .\control_reg[3] (control_reg_adj_916[3]), 
            .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), 
            .\read_size[2] (read_size_adj_920[2]), .n29768(n29768), .\steps_reg[9] (steps_reg_adj_918[9]), 
            .\steps_reg[6] (steps_reg_adj_918[6]), .\steps_reg[5] (steps_reg_adj_918[5]), 
            .\steps_reg[3] (steps_reg_adj_918[3]), .n32(n32_adj_542), .n29770(n29770), 
            .read_value({read_value_adj_919}), .n4071(n4071), .limit_c_1(limit_c_1), 
            .n8476(n8475[7]), .n29788(n29788), .n31921(n31921), .n21084(n21084), 
            .n21092(n21092), .n6785(n6756[3]), .int_step(int_step), .n22(n22), 
            .n31919(n31919), .n31905(n31905), .n16545(n16545), .n7996(n7996), 
            .n8030(n8030)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(599[25] 612[45])
    LUT4 m1_lut (.Z(n33682)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.read_value({read_value_adj_1001}), 
            .debug_c_c(debug_c_c), .n2850(n2850), .n31991(n31991), .n3899({n3899}), 
            .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_1002[0]), .n29798(n29798), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .n22330(n22330), .n579(n571_adj_1020[0]), .limit_latched(limit_latched_adj_683), 
            .prev_limit_latched(prev_limit_latched_adj_684), .n14661(n14661), 
            .prev_select(prev_select_adj_719), .n31938(n31938), .n32(n32), 
            .n32_adj_37(n32_adj_543), .prev_step_clk(prev_step_clk_adj_637), 
            .step_clk(step_clk_adj_636), .n31918(n31918), .n22(n22_adj_585), 
            .n32_adj_38(n32_adj_542), .prev_step_clk_adj_39(prev_step_clk_adj_590), 
            .step_clk_adj_40(step_clk_adj_589), .n31919(n31919), .n22_adj_41(n22), 
            .prev_step_clk_adj_42(prev_step_clk), .n34(n34), .step_clk_adj_43(step_clk), 
            .n31920(n31920), .n24(n24), .\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .\read_size[2] (read_size_adj_1002[2]), 
            .n94(n94_adj_819), .Stepper_A_M1_c_1(Stepper_A_M1_c_1), .n13710(n13710), 
            .\databus[1] (databus[1]), .Stepper_A_M2_c_2(Stepper_A_M2_c_2), 
            .\databus[2] (databus[2]), .\databus[3] (databus[3]), .\databus[4] (databus[4]), 
            .Stepper_A_Dir_c(Stepper_A_Dir_c), .\databus[5] (databus[5]), 
            .Stepper_A_En_c(Stepper_A_En_c), .\databus[6] (databus[6]), 
            .\control_reg[7] (control_reg_adj_998[7]), .n11981(n11981), 
            .\databus[7] (databus[7]), .n31910(n31910), .\databus[8] (databus[8]), 
            .\databus[9] (databus[9]), .\databus[10] (databus[10]), .\databus[11] (databus[11]), 
            .\databus[12] (databus[12]), .\databus[13] (databus[13]), .\databus[14] (databus[14]), 
            .\databus[15] (databus[15]), .\databus[16] (databus[16]), .\databus[17] (databus[17]), 
            .\databus[18] (databus[18]), .\databus[19] (databus[19]), .\databus[20] (databus[20]), 
            .\databus[21] (databus[21]), .\databus[22] (databus[22]), .\databus[23] (databus[23]), 
            .\databus[24] (databus[24]), .\databus[25] (databus[25]), .\databus[26] (databus[26]), 
            .\databus[27] (databus[27]), .\databus[28] (databus[28]), .\databus[29] (databus[29]), 
            .\databus[30] (databus[30]), .\databus[31] (databus[31]), .n224({n224_adj_1006}), 
            .n31911(n31911), .n32056(n32056), .n13323(n13323), .n32003(n32003), 
            .n30489(n30489), .limit_c_3(limit_c_3), .n27766(n27766), .Stepper_A_Step_c(Stepper_A_Step_c), 
            .n8494(n8493[7]), .n31903(n31903), .n16566(n16566), .n8204(n8204), 
            .n8238(n8238)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(629[25] 642[45])
    LUT4 i6_2_lut (.A(state_adj_1082[1]), .B(state_adj_1082[0]), .Z(n7645[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    defparam i6_2_lut.init = 16'h6666;
    ClockDivider_U10 pwm_clk_div (.GND_net(GND_net), .clk_255kHz(clk_255kHz), 
            .debug_c_c(debug_c_c), .n241(n241), .n31991(n31991), .n7718(n7718), 
            .n30378(n30378), .n14374(n14374), .n30518(n30518), .n27956(n27956), 
            .n30516(n30516), .n27960(n27960), .n30381(n30381), .n13735(n13735), 
            .n30505(n30505), .n14315(n14315), .n30445(n30445), .n14358(n14358), 
            .n30514(n30514), .n27757(n27757), .n2816(n2816), .n7753(n7753), 
            .n30426(n30426), .n14369(n14369), .n30510(n30510), .n27759(n27759), 
            .n30520(n30520), .n27883(n27883), .n30512(n30512), .n27758(n27758)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(544[15] 547[41])
    LUT4 i1_2_lut_rep_292 (.A(n8343), .B(select_clk), .Z(n31909)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(471[17:42])
    defparam i1_2_lut_rep_292.init = 16'h2222;
    LUT4 i20_2_lut_rep_307_3_lut_4_lut (.A(n32003), .B(n13323), .C(n33683), 
         .D(select[4]), .Z(n31924)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(552[4] 581[11])
    defparam i20_2_lut_rep_307_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_3_lut_rep_290_4_lut (.A(n8343), .B(select_clk), .C(state_adj_1082[0]), 
         .D(n31991), .Z(n31907)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(471[17:42])
    defparam i1_3_lut_rep_290_4_lut.init = 16'h0002;
    LUT4 i23204_4_lut_4_lut (.A(n1153), .B(n1165), .C(n29869), .D(n31948), 
         .Z(n30516)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+!(D))) */ ;
    defparam i23204_4_lut_4_lut.init = 16'hbb02;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n31991), .B(prev_select_adj_719), 
         .C(n31970), .D(select[4]), .Z(n2850)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    \ClockDividerP_SP(factor=120000)  clk_100Hz_divider (.debug_c_0(debug_c_0), 
            .debug_c_c(debug_c_c), .n31991(n31991), .n2853(n2853), .n30361(n30361), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(647[29] 649[61])
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.read_value({read_value_adj_960}), 
            .debug_c_c(debug_c_c), .n13876(n13876), .GND_net(GND_net), 
            .VCC_net(VCC_net), .Stepper_Z_nFault_c(Stepper_Z_nFault_c), 
            .\read_size[0] (read_size_adj_961[0]), .n29175(n29175), .n31991(n31991), 
            .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n110(n110), .n579(n571_adj_1020[0]), 
            .prev_step_clk(prev_step_clk_adj_637), .step_clk(step_clk_adj_636), 
            .limit_latched(limit_latched_adj_634), .prev_limit_latched(prev_limit_latched_adj_635), 
            .n13698(n13698), .prev_select(prev_select_adj_672), .n31982(n31982), 
            .databus({databus}), .n3984(n3984), .\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .n27787(n27787), .\read_size[2] (read_size_adj_961[2]), 
            .n29174(n29174), .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), .n13693(n13693), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .Stepper_Z_Dir_c(Stepper_Z_Dir_c), 
            .Stepper_Z_En_c(Stepper_Z_En_c), .\control_reg[7] (control_reg_adj_957[7]), 
            .n11020(n11020), .n9139(n9139), .n32(n32_adj_543), .n22(n22_adj_585), 
            .n31918(n31918), .limit_c_2(limit_c_2), .Stepper_Z_Step_c(Stepper_Z_Step_c), 
            .n8485(n8484[7]), .n8100(n8100), .n31902(n31902), .n16565(n16565), 
            .n8134(n8134)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(614[25] 627[45])
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.\read_size[2] (read_size_adj_908[2]), 
            .debug_c_c(debug_c_c), .n13708(n13708), .n31933(n31933), .databus({databus}), 
            .n4168(n4168), .n31991(n31991), .\register_addr[0] (register_addr[0]), 
            .n13647(n13647), .\read_size[0] (read_size_adj_908[0]), .n31922(n31922), 
            .Stepper_X_M0_c_0(Stepper_X_M0_c_0), .n14258(n14258), .n579(n571_adj_1020[0]), 
            .prev_step_clk(prev_step_clk), .step_clk(step_clk), .limit_latched(limit_latched), 
            .prev_limit_latched(prev_limit_latched), .prev_select(prev_select_adj_583), 
            .n31951(n31951), .Stepper_X_Step_c(Stepper_X_Step_c), .n27768(n27768), 
            .\register_addr[1] (register_addr[1]), .GND_net(GND_net), .n34(n34), 
            .n31915(n31915), .n608(n580[4]), .n610(n580[2]), .n1(n1), 
            .\control_reg[7] (control_reg[7]), .n13642(n13642), .n10962(n10962), 
            .Stepper_X_En_c(Stepper_X_En_c), .Stepper_X_Dir_c(Stepper_X_Dir_c), 
            .Stepper_X_M2_c_2(Stepper_X_M2_c_2), .Stepper_X_M1_c_1(Stepper_X_M1_c_1), 
            .read_value({read_value_adj_907}), .VCC_net(VCC_net), .Stepper_X_nFault_c(Stepper_X_nFault_c), 
            .limit_c_0(limit_c_0), .n24(n24), .n31920(n31920), .n31904(n31904), 
            .n16744(n16744), .n7892(n7892), .n7926(n7926)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(584[25] 597[45])
    EncoderPeripheral right_encoder (.\read_size[0] (read_size_adj_1049[0]), 
            .debug_c_c(debug_c_c), .n14116(n14116), .n31950(n31950), .n31986(n31986), 
            .prev_select(prev_select_adj_797), .n31990(n31990), .read_value({read_value_adj_1048}), 
            .\register_addr[0] (register_addr[0]), .\read_size[2] (read_size_adj_1049[2]), 
            .n5(n9_adj_1320[1]), .encoder_ra_c(encoder_ra_c), .encoder_rb_c(encoder_rb_c), 
            .encoder_ri_c(encoder_ri_c), .n13779(n13779), .n97(n99_adj_1308[0]), 
            .\quadB_delayed[2] (quadB_delayed_adj_1139[2]), .\quadA_delayed[1] (quadA_delayed_adj_1138[1]), 
            .GND_net(GND_net), .n31952(n31952), .n4433(n4401[0]), .VCC_net(VCC_net), 
            .\quadB_delayed[1] (quadB_delayed_adj_1139[1]), .\quadA_delayed[2] (quadA_delayed_adj_1138[2])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(686[20] 696[47])
    \ProtocolInterface(baud_div=12)  protocol_interface (.databus({databus}), 
            .register_addr({Open_7, Open_8, register_addr[5:0]}), .n32090(n32090), 
            .n30166(n30166), .debug_c_c(debug_c_c), .\select[7] (select[7]), 
            .n31975(n31975), .n32001(n32001), .prev_select(prev_select_adj_760), 
            .n31923(n31923), .\select[4] (select[4]), .\select[3] (select[3]), 
            .\select[2] (select[2]), .\select[1] (select[1]), .databus_out({databus_out}), 
            .n13608(n13608), .n32075(n32075), .rw(rw), .n31926(n31926), 
            .n1486(n1468[14]), .debug_c_7(debug_c_7), .n31928(n31928), 
            .n31911(n31911), .n224({n224_adj_1006}), .n3899({n3899}), 
            .prev_select_adj_1(prev_select_adj_672), .n31991(n31991), .n13876(n13876), 
            .\sendcount[1] (sendcount[1]), .n32052(n32052), .n8(n8_adj_584), 
            .n31944(n31944), .n32032(n32032), .n32089(n32089), .n29768(n29768), 
            .n32011(n32011), .n29174(n29174), .n29175(n29175), .n31996(n31996), 
            .n31965(n31965), .\read_value[1] (read_value_adj_907[1]), .n4(n4), 
            .n13700(n13700), .n31972(n31972), .n29770(n29770), .n32056(n32056), 
            .n11158(n11158), .prev_select_adj_2(prev_select_adj_625), .n31986(n31986), 
            .\read_value[28] (read_value_adj_919[28]), .n33683(n33683), 
            .n3(n3_adj_626), .n27768(n27768), .\control_reg[7] (control_reg[7]), 
            .n32088(n32088), .n34(n34), .n31933(n31933), .n29916(n29916), 
            .n13647(n13647), .n32005(n32005), .\register[2][3] (\register[2] [3]), 
            .n5980(n5951[3]), .n27787(n27787), .\control_reg[7]_adj_3 (control_reg_adj_957[7]), 
            .n32(n32_adj_543), .prev_select_adj_4(prev_select_adj_583), 
            .n27886(n27886), .n33682(n33682), .n13323(n13323), .n31938(n31938), 
            .\read_value[27] (read_value_adj_919[27]), .n3_adj_5(n3_adj_821), 
            .n29798(n29798), .n31937(n31937), .n33680(n33680), .n15(n15_adj_855), 
            .n31940(n31940), .n250_adj_6(n250), .n32034(n32034), .n31982(n31982), 
            .n31955(n31955), .n4071(n4071), .n13708(n13708), .n32003(n32003), 
            .n94(n94_adj_819), .n32006(n32006), .\register[2][4] (\register[2] [4]), 
            .n29197(n29197), .\register[2][5] (\register[2] [5]), .n29211(n29211), 
            .\register[2][6] (\register[2] [6]), .n29213(n29213), .\register[2][7] (\register[2] [7]), 
            .n29207(n29207), .\register[2][8] (\register[2] [8]), .n29199(n29199), 
            .\register[2][9] (\register[2] [9]), .n29215(n29215), .\register[2][10] (\register[2] [10]), 
            .n29189(n29189), .n31915(n31915), .n31990(n31990), .\register[2][11] (\register[2] [11]), 
            .n29190(n29190), .\register[2][12] (\register[2] [12]), .n29201(n29201), 
            .\register[2][13] (\register[2] [13]), .n29209(n29209), .\register[2][14] (\register[2] [14]), 
            .n29203(n29203), .n14372(n14372), .n9362(n9362), .n12930(n12930), 
            .\register[2][15] (\register[2] [15]), .n29191(n29191), .\register[2][16] (\register[2] [16]), 
            .n29193(n29193), .n22(n22_adj_631), .n12(n12_adj_847), .n8_adj_7(n8_adj_848), 
            .\register[2][17] (\register[2] [17]), .n29205(n29205), .\reg_size[2] (reg_size[2]), 
            .n32068(n32068), .n32004(n32004), .n5811(n5811), .n27946(n27946), 
            .n31951(n31951), .n52(n52), .\register[2][18] (\register[2] [18]), 
            .n29194(n29194), .n1480(n1468[20]), .n31977(n31977), .\register[2][19] (\register[2] [19]), 
            .n29196(n29196), .\register[2][20] (\register[2] [20]), .n29198(n29198), 
            .\register[2][21] (\register[2] [21]), .n29200(n29200), .n1483(n1468[17]), 
            .\register[2][22] (\register[2] [22]), .n29202(n29202), .\register[2][23] (\register[2] [23]), 
            .n29204(n29204), .n32030(n32030), .\register[2][24] (\register[2] [24]), 
            .n29206(n29206), .\register[2][25] (\register[2] [25]), .n29208(n29208), 
            .\register[2][26] (\register[2] [26]), .n29210(n29210), .\register[2][27] (\register[2] [27]), 
            .n29214(n29214), .n4_adj_8(n4_adj_833), .\register[2][28] (\register[2] [28]), 
            .n29216(n29216), .\register[2][29] (\register[2] [29]), .n29195(n29195), 
            .\register[2][30] (\register[2] [30]), .n29192(n29192), .\register[2][31] (\register[2] [31]), 
            .n29212(n29212), .n31987(n31987), .n31953(n31953), .n14094(n14094), 
            .n31970(n31970), .n31910(n31910), .n13710(n13710), .\read_value[26] (read_value_adj_919[26]), 
            .n3_adj_9(n3_adj_817), .\read_value[25] (read_value_adj_919[25]), 
            .n3_adj_10(n3_adj_677), .\read_value[24] (read_value_adj_919[24]), 
            .n3_adj_11(n3_adj_814), .\steps_reg[5] (steps_reg_adj_918[5]), 
            .n14(n14), .\steps_reg[6] (steps_reg_adj_918[6]), .n13(n13), 
            .\steps_reg[3] (steps_reg_adj_918[3]), .n12_adj_12(n12), .\read_value[23] (read_value_adj_919[23]), 
            .n3_adj_13(n3_adj_803), .\read_value[22] (read_value_adj_919[22]), 
            .n3_adj_14(n3_adj_676), .\control_reg[7]_adj_15 (control_reg_adj_998[7]), 
            .n8494(n8493[7]), .\read_value[21] (read_value_adj_919[21]), 
            .n3_adj_16(n3_adj_824), .\read_value[20] (read_value_adj_919[20]), 
            .n3_adj_17(n3_adj_673), .\read_value[19] (read_value_adj_919[19]), 
            .n3_adj_18(n3_adj_761), .\read_value[18] (read_value_adj_919[18]), 
            .n3_adj_19(n3_adj_674), .n13642(n13642), .\control_reg[7]_adj_20 (control_reg_adj_916[7]), 
            .n8476(n8475[7]), .\read_value[17] (read_value_adj_919[17]), 
            .n3_adj_21(n3_adj_629), .\read_value[16] (read_value_adj_919[16]), 
            .n3_adj_22(n3_adj_628), .\read_value[15] (read_value_adj_919[15]), 
            .n3_adj_23(n3_adj_856), .\read_value[14] (read_value_adj_919[14]), 
            .n3_adj_24(n3), .n13667(n13667), .\read_value[13] (read_value_adj_919[13]), 
            .n3_adj_25(n3_adj_862), .n3984(n3984), .\read_value[12] (read_value_adj_919[12]), 
            .n3_adj_26(n3_adj_825), .\read_value[11] (read_value_adj_919[11]), 
            .n3_adj_27(n3_adj_827), .n13693(n13693), .n9139(n9139), .n1(n1), 
            .n31942(n31942), .\read_value[10] (read_value_adj_919[10]), 
            .n3_adj_28(n3_adj_838), .\read_value[9] (read_value_adj_919[9]), 
            .n3_adj_29(n3_adj_840), .\read_value[8] (read_value_adj_919[8]), 
            .n3_adj_30(n3_adj_829), .debug_c_2(debug_c_2), .debug_c_3(debug_c_3), 
            .n27766(n27766), .n32_adj_31(n32), .debug_c_4(debug_c_4), 
            .debug_c_5(debug_c_5), .n31921(n31921), .n14661(n14661), .n31922(n31922), 
            .n96(n96_adj_823), .\read_value[31] (read_value_adj_919[31]), 
            .n3_adj_32(n3_adj_805), .\read_value[29] (read_value_adj_919[29]), 
            .n3_adj_33(n3_adj_801), .n8485(n8484[7]), .\read_value[30] (read_value_adj_919[30]), 
            .n3_adj_34(n3_adj_799), .prev_select_adj_35(prev_select_adj_797), 
            .n5(n9_adj_1320[1]), .n27769(n27769), .n32_adj_36(n32_adj_542), 
            .\reset_count[14] (reset_count[14]), .\reset_count[13] (reset_count[13]), 
            .\reset_count[12] (reset_count[12]), .n29900(n29900), .n10889(n10889), 
            .GND_net(GND_net), .uart_rx_c(uart_rx_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(499[26] 509[57])
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (debug_c_c, n9312, n31991, read_size, 
            n14372, n27946, \register[2][31] , \register[2][30] , \register[2][29] , 
            prev_clk_1Hz, clk_1Hz, \register[2][28] , \register[2][27] , 
            prev_select, \select[1] , \register[2][26] , \register[2][25] , 
            \register[2][24] , \register[2][23] , \register[2][22] , \register[2][21] , 
            \register[2][20] , \register[2][19] , \register[2][18] , \register[2][17] , 
            \register[2][16] , \register[2][15] , \register[2][14] , \register[2][13] , 
            \register[2][12] , \register[2][11] , \register[2][10] , \register[2][9] , 
            \register[2][8] , \register[2][7] , \register[2][6] , \register[2][5] , 
            \register[2][4] , \register[2][3] , rw, n46, n11158, \register_addr[1] , 
            \register_addr[0] , n32034, \register_addr[5] , n32032, 
            \databus[1] , timeout_pause, n32088, signal_light_c, \register[0][7] , 
            n32016, n8, n31937, read_value, n9362, GND_net, xbee_pause_c, 
            n5980, n29197, n29211, n29213, n29207, n29199, n29215, 
            n29189, n29190, n29201, n29209, n29203, n29191, n29193, 
            n29205, n29194, n29196, n29198, n29200, n29202, n29204, 
            n29206, n29208, n29210, n250, n15, n29214, n29216, 
            n29195, n29192, n31965, n31975, n29212, n32052, n32005, 
            n31972, n2863, n30358) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n9312;
    input n31991;
    output [2:0]read_size;
    input n14372;
    input n27946;
    output \register[2][31] ;
    output \register[2][30] ;
    output \register[2][29] ;
    output prev_clk_1Hz;
    output clk_1Hz;
    output \register[2][28] ;
    output \register[2][27] ;
    output prev_select;
    input \select[1] ;
    output \register[2][26] ;
    output \register[2][25] ;
    output \register[2][24] ;
    output \register[2][23] ;
    output \register[2][22] ;
    output \register[2][21] ;
    output \register[2][20] ;
    output \register[2][19] ;
    output \register[2][18] ;
    output \register[2][17] ;
    output \register[2][16] ;
    output \register[2][15] ;
    output \register[2][14] ;
    output \register[2][13] ;
    output \register[2][12] ;
    output \register[2][11] ;
    output \register[2][10] ;
    output \register[2][9] ;
    output \register[2][8] ;
    output \register[2][7] ;
    output \register[2][6] ;
    output \register[2][5] ;
    output \register[2][4] ;
    output \register[2][3] ;
    input rw;
    output n46;
    input n11158;
    input \register_addr[1] ;
    input \register_addr[0] ;
    input n32034;
    input \register_addr[5] ;
    input n32032;
    input \databus[1] ;
    input timeout_pause;
    output n32088;
    output signal_light_c;
    input \register[0][7] ;
    output n32016;
    input n8;
    input n31937;
    output [31:0]read_value;
    input n9362;
    input GND_net;
    input xbee_pause_c;
    input n5980;
    input n29197;
    input n29211;
    input n29213;
    input n29207;
    input n29199;
    input n29215;
    input n29189;
    input n29190;
    input n29201;
    input n29209;
    input n29203;
    input n29191;
    input n29193;
    input n29205;
    input n29194;
    input n29196;
    input n29198;
    input n29200;
    input n29202;
    input n29204;
    input n29206;
    input n29208;
    input n29210;
    input n250;
    input n15;
    input n29214;
    input n29216;
    input n29195;
    input n29192;
    input n31965;
    input n31975;
    input n29212;
    input n32052;
    input n32005;
    input n31972;
    input n2863;
    output n30358;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    wire [31:0]n100;
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    
    wire n179, n1, n2;
    wire [31:0]n100_adj_540;
    
    wire force_pause, n31897, n31898, n28580, n27021, n27020, n27019, 
        n27018, n27017, n27016, n27015, n27014, n27013, n27012, 
        n27011, n27010, n27009, n27008, n27007, n27006, n27548, 
        n16493;
    wire [31:0]n5951;
    
    wire n11160;
    
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n27946), .SP(n14372), .CK(debug_c_c), 
            .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][31] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][30] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][29] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_150 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam prev_clk_1Hz_150.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_151 (.D(n179), .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam xbee_pause_latched_151.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][28] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][27] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1S3AX prev_select_149 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam prev_select_149.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][26] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][25] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][23] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][22] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][21] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][19] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][18] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][17] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n9312), .CD(n31991), 
            .CK(debug_c_c), .Q(\register[2][10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2][9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2][8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2][7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2][6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2][5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2][3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n9312), .CD(n31991), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    LUT4 i14_2_lut (.A(\select[1] ), .B(rw), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(36[19:32])
    defparam i14_2_lut.init = 16'h8888;
    LUT4 i14979_4_lut (.A(n1), .B(n11158), .C(n2), .D(\register_addr[1] ), 
         .Z(n100_adj_540[1])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i14979_4_lut.init = 16'h3022;
    LUT4 i15063_2_lut (.A(force_pause), .B(\register_addr[0] ), .Z(n1)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15063_2_lut.init = 16'heeee;
    LUT4 i15315_2_lut (.A(\register[2] [1]), .B(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i15315_2_lut.init = 16'h2222;
    LUT4 register_addr_0__bdd_4_lut_24345 (.A(\register_addr[0] ), .B(\register[0] [2]), 
         .C(\register_addr[1] ), .D(\register[2] [2]), .Z(n31897)) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam register_addr_0__bdd_4_lut_24345.init = 16'h5e0e;
    LUT4 n31897_bdd_2_lut_4_lut (.A(n32034), .B(\register_addr[5] ), .C(n32032), 
         .D(n31897), .Z(n31898)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam n31897_bdd_2_lut_4_lut.init = 16'h0100;
    FD1P3IX force_pause_152 (.D(\databus[1] ), .SP(n28580), .CD(n31991), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam force_pause_152.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_471 (.A(timeout_pause), .B(force_pause), .C(\register[0] [2]), 
         .Z(n32088)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(39[24:72])
    defparam i2_3_lut_rep_471.init = 16'hfefe;
    LUT4 i14672_2_lut_4_lut (.A(timeout_pause), .B(force_pause), .C(\register[0] [2]), 
         .D(clk_1Hz), .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(39[24:72])
    defparam i14672_2_lut_4_lut.init = 16'hfffe;
    LUT4 i15151_2_lut_rep_399_4_lut (.A(timeout_pause), .B(force_pause), 
         .C(\register[0] [2]), .D(\register[0][7] ), .Z(n32016)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(39[24:72])
    defparam i15151_2_lut_rep_399_4_lut.init = 16'h0100;
    LUT4 i1_4_lut (.A(prev_select), .B(n31991), .C(n8), .D(n31937), 
         .Z(n28580)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'hccdc;
    FD1P3AX read_value__i2 (.D(n31898), .SP(n14372), .CK(debug_c_c), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n100_adj_540[1]), .SP(n14372), .CD(n9362), 
            .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i1.GSR = "ENABLED";
    CCU2D add_135_33 (.A0(\register[2][31] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27021), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_33.INIT0 = 16'h5aaa;
    defparam add_135_33.INIT1 = 16'h0000;
    defparam add_135_33.INJECT1_0 = "NO";
    defparam add_135_33.INJECT1_1 = "NO";
    CCU2D add_135_31 (.A0(\register[2][29] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][30] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27020), .COUT(n27021), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_31.INIT0 = 16'h5aaa;
    defparam add_135_31.INIT1 = 16'h5aaa;
    defparam add_135_31.INJECT1_0 = "NO";
    defparam add_135_31.INJECT1_1 = "NO";
    CCU2D add_135_29 (.A0(\register[2][27] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][28] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27019), .COUT(n27020), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_29.INIT0 = 16'h5aaa;
    defparam add_135_29.INIT1 = 16'h5aaa;
    defparam add_135_29.INJECT1_0 = "NO";
    defparam add_135_29.INJECT1_1 = "NO";
    CCU2D add_135_27 (.A0(\register[2][25] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][26] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27018), .COUT(n27019), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_27.INIT0 = 16'h5aaa;
    defparam add_135_27.INIT1 = 16'h5aaa;
    defparam add_135_27.INJECT1_0 = "NO";
    defparam add_135_27.INJECT1_1 = "NO";
    CCU2D add_135_25 (.A0(\register[2][23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27017), .COUT(n27018), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_25.INIT0 = 16'h5aaa;
    defparam add_135_25.INIT1 = 16'h5aaa;
    defparam add_135_25.INJECT1_0 = "NO";
    defparam add_135_25.INJECT1_1 = "NO";
    CCU2D add_135_23 (.A0(\register[2][21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27016), .COUT(n27017), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_23.INIT0 = 16'h5aaa;
    defparam add_135_23.INIT1 = 16'h5aaa;
    defparam add_135_23.INJECT1_0 = "NO";
    defparam add_135_23.INJECT1_1 = "NO";
    CCU2D add_135_21 (.A0(\register[2][19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27015), .COUT(n27016), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_21.INIT0 = 16'h5aaa;
    defparam add_135_21.INIT1 = 16'h5aaa;
    defparam add_135_21.INJECT1_0 = "NO";
    defparam add_135_21.INJECT1_1 = "NO";
    CCU2D add_135_19 (.A0(\register[2][17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27014), .COUT(n27015), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_19.INIT0 = 16'h5aaa;
    defparam add_135_19.INIT1 = 16'h5aaa;
    defparam add_135_19.INJECT1_0 = "NO";
    defparam add_135_19.INJECT1_1 = "NO";
    CCU2D add_135_17 (.A0(\register[2][15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27013), .COUT(n27014), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_17.INIT0 = 16'h5aaa;
    defparam add_135_17.INIT1 = 16'h5aaa;
    defparam add_135_17.INJECT1_0 = "NO";
    defparam add_135_17.INJECT1_1 = "NO";
    CCU2D add_135_15 (.A0(\register[2][13] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][14] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27012), .COUT(n27013), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_15.INIT0 = 16'h5aaa;
    defparam add_135_15.INIT1 = 16'h5aaa;
    defparam add_135_15.INJECT1_0 = "NO";
    defparam add_135_15.INJECT1_1 = "NO";
    CCU2D add_135_13 (.A0(\register[2][11] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][12] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27011), .COUT(n27012), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_13.INIT0 = 16'h5aaa;
    defparam add_135_13.INIT1 = 16'h5aaa;
    defparam add_135_13.INJECT1_0 = "NO";
    defparam add_135_13.INJECT1_1 = "NO";
    CCU2D add_135_11 (.A0(\register[2][9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][10] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27010), .COUT(n27011), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_11.INIT0 = 16'h5aaa;
    defparam add_135_11.INIT1 = 16'h5aaa;
    defparam add_135_11.INJECT1_0 = "NO";
    defparam add_135_11.INJECT1_1 = "NO";
    CCU2D add_135_9 (.A0(\register[2][7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][8] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27009), .COUT(n27010), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_9.INIT0 = 16'h5aaa;
    defparam add_135_9.INIT1 = 16'h5aaa;
    defparam add_135_9.INJECT1_0 = "NO";
    defparam add_135_9.INJECT1_1 = "NO";
    CCU2D add_135_7 (.A0(\register[2][5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27008), .COUT(n27009), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_7.INIT0 = 16'h5aaa;
    defparam add_135_7.INIT1 = 16'h5aaa;
    defparam add_135_7.INJECT1_0 = "NO";
    defparam add_135_7.INJECT1_1 = "NO";
    CCU2D add_135_5 (.A0(\register[2][3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27007), .COUT(n27008), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_5.INIT0 = 16'h5aaa;
    defparam add_135_5.INIT1 = 16'h5aaa;
    defparam add_135_5.INJECT1_0 = "NO";
    defparam add_135_5.INJECT1_1 = "NO";
    CCU2D add_135_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27006), .COUT(n27007), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_3.INIT0 = 16'h5aaa;
    defparam add_135_3.INIT1 = 16'h5aaa;
    defparam add_135_3.INJECT1_0 = "NO";
    defparam add_135_3.INJECT1_1 = "NO";
    LUT4 i115_1_lut (.A(xbee_pause_c), .Z(n179)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(55[26:39])
    defparam i115_1_lut.init = 16'h5555;
    CCU2D add_135_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27006), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(104[23:39])
    defparam add_135_1.INIT0 = 16'hF000;
    defparam add_135_1.INIT1 = 16'h5555;
    defparam add_135_1.INJECT1_0 = "NO";
    defparam add_135_1.INJECT1_1 = "NO";
    FD1P3IX read_value__i3 (.D(n5980), .SP(n14372), .CD(n9362), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29197), .SP(n14372), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29211), .SP(n14372), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29213), .SP(n14372), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29207), .SP(n14372), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29199), .SP(n14372), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29215), .SP(n14372), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29189), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29190), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29201), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29209), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29203), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29191), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29193), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29205), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29194), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29196), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29198), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29200), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29202), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29204), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29206), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29208), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29210), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_size_i0_i1 (.D(n250), .SP(n14372), .CD(n27548), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n15), .SP(n14372), .CD(n16493), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29214), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29216), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29195), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29192), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n5951[0]), .SP(n14372), .CD(n9362), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(\register_addr[0] ), .B(n14372), .C(\register_addr[1] ), 
         .D(n31965), .Z(n27548)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!B))) */ ;
    defparam i2_4_lut.init = 16'h00c4;
    LUT4 i9862_4_lut (.A(n14372), .B(\register_addr[0] ), .C(n31975), 
         .D(\register_addr[1] ), .Z(n16493)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;
    defparam i9862_4_lut.init = 16'ha0a8;
    FD1P3AX read_value__i31 (.D(n29212), .SP(n14372), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=520, LSE_RLINE=531 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(51[9] 106[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i14621_4_lut (.A(n32052), .B(n32005), .C(n11160), .D(n31972), 
         .Z(n5951[0])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;
    defparam i14621_4_lut.init = 16'hccdc;
    LUT4 i4534_3_lut (.A(n32088), .B(\register[2] [0]), .C(\register_addr[1] ), 
         .Z(n11160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4534_3_lut.init = 16'hcaca;
    \ClockDividerP(factor=12000000)  uptime_div (.clk_1Hz(clk_1Hz), .debug_c_c(debug_c_c), 
            .n31991(n31991), .n2863(n2863), .n30358(n30358), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(108[28] 110[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (clk_1Hz, debug_c_c, n31991, n2863, 
            n30358, GND_net) /* synthesis syn_module_defined=1 */ ;
    output clk_1Hz;
    input debug_c_c;
    input n31991;
    input n2863;
    output n30358;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n7822;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n27, n27734, n25, n26, n24, n19, n32, n28, n20, n29, 
        n26_adj_537, n27347, n27346, n27345, n27344, n27343, n27342, 
        n27341, n27340, n27339, n27338, n27337, n27336, n27335, 
        n27334, n27333, n27332, n27507, n27506, n27505, n27504, 
        n27503, n27502, n27501, n27500, n27499, n27498, n27497, 
        n27496;
    
    FD1S3IX clk_o_14 (.D(n7822), .CK(debug_c_c), .CD(n31991), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2635__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2863), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i0.GSR = "ENABLED";
    LUT4 i23046_4_lut (.A(n27), .B(n27734), .C(n25), .D(n26), .Z(n30358)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i23046_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n27734)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_537), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_472 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_472.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_473 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_473.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_537)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    CCU2D count_2635_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27347), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_33.INIT1 = 16'h0000;
    defparam count_2635_add_4_33.INJECT1_0 = "NO";
    defparam count_2635_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27346), .COUT(n27347), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_31.INJECT1_0 = "NO";
    defparam count_2635_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27345), .COUT(n27346), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_29.INJECT1_0 = "NO";
    defparam count_2635_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27344), .COUT(n27345), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_27.INJECT1_0 = "NO";
    defparam count_2635_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27343), .COUT(n27344), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_25.INJECT1_0 = "NO";
    defparam count_2635_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27342), .COUT(n27343), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_23.INJECT1_0 = "NO";
    defparam count_2635_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27341), .COUT(n27342), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_21.INJECT1_0 = "NO";
    defparam count_2635_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27340), .COUT(n27341), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_19.INJECT1_0 = "NO";
    defparam count_2635_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27339), .COUT(n27340), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_17.INJECT1_0 = "NO";
    defparam count_2635_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27338), .COUT(n27339), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_15.INJECT1_0 = "NO";
    defparam count_2635_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27337), .COUT(n27338), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_13.INJECT1_0 = "NO";
    defparam count_2635_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27336), .COUT(n27337), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_11.INJECT1_0 = "NO";
    defparam count_2635_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27335), .COUT(n27336), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_9.INJECT1_0 = "NO";
    defparam count_2635_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27334), .COUT(n27335), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_7.INJECT1_0 = "NO";
    defparam count_2635_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27333), .COUT(n27334), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_5.INJECT1_0 = "NO";
    defparam count_2635_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27332), .COUT(n27333), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2635_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2635_add_4_3.INJECT1_0 = "NO";
    defparam count_2635_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2635_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27332), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635_add_4_1.INIT0 = 16'hF000;
    defparam count_2635_add_4_1.INIT1 = 16'h0555;
    defparam count_2635_add_4_1.INJECT1_0 = "NO";
    defparam count_2635_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2635__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2863), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i1.GSR = "ENABLED";
    FD1S3IX count_2635__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2863), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i2.GSR = "ENABLED";
    FD1S3IX count_2635__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2863), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i3.GSR = "ENABLED";
    FD1S3IX count_2635__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2863), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i4.GSR = "ENABLED";
    FD1S3IX count_2635__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2863), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i5.GSR = "ENABLED";
    FD1S3IX count_2635__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2863), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i6.GSR = "ENABLED";
    FD1S3IX count_2635__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2863), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i7.GSR = "ENABLED";
    FD1S3IX count_2635__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2863), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i8.GSR = "ENABLED";
    FD1S3IX count_2635__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2863), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i9.GSR = "ENABLED";
    FD1S3IX count_2635__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i10.GSR = "ENABLED";
    FD1S3IX count_2635__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i11.GSR = "ENABLED";
    FD1S3IX count_2635__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i12.GSR = "ENABLED";
    FD1S3IX count_2635__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i13.GSR = "ENABLED";
    FD1S3IX count_2635__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i14.GSR = "ENABLED";
    FD1S3IX count_2635__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i15.GSR = "ENABLED";
    FD1S3IX count_2635__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i16.GSR = "ENABLED";
    FD1S3IX count_2635__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i17.GSR = "ENABLED";
    FD1S3IX count_2635__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i18.GSR = "ENABLED";
    FD1S3IX count_2635__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i19.GSR = "ENABLED";
    FD1S3IX count_2635__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i20.GSR = "ENABLED";
    FD1S3IX count_2635__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i21.GSR = "ENABLED";
    FD1S3IX count_2635__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i22.GSR = "ENABLED";
    FD1S3IX count_2635__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i23.GSR = "ENABLED";
    FD1S3IX count_2635__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i24.GSR = "ENABLED";
    FD1S3IX count_2635__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i25.GSR = "ENABLED";
    FD1S3IX count_2635__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i26.GSR = "ENABLED";
    FD1S3IX count_2635__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i27.GSR = "ENABLED";
    FD1S3IX count_2635__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i28.GSR = "ENABLED";
    FD1S3IX count_2635__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i29.GSR = "ENABLED";
    FD1S3IX count_2635__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i30.GSR = "ENABLED";
    FD1S3IX count_2635__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2863), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2635__i31.GSR = "ENABLED";
    CCU2D add_20099_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27507), 
          .S0(n7822));
    defparam add_20099_cout.INIT0 = 16'h0000;
    defparam add_20099_cout.INIT1 = 16'h0000;
    defparam add_20099_cout.INJECT1_0 = "NO";
    defparam add_20099_cout.INJECT1_1 = "NO";
    CCU2D add_20099_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27506), .COUT(n27507));
    defparam add_20099_24.INIT0 = 16'h5555;
    defparam add_20099_24.INIT1 = 16'h5555;
    defparam add_20099_24.INJECT1_0 = "NO";
    defparam add_20099_24.INJECT1_1 = "NO";
    CCU2D add_20099_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27505), .COUT(n27506));
    defparam add_20099_22.INIT0 = 16'h5555;
    defparam add_20099_22.INIT1 = 16'h5555;
    defparam add_20099_22.INJECT1_0 = "NO";
    defparam add_20099_22.INJECT1_1 = "NO";
    CCU2D add_20099_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27504), .COUT(n27505));
    defparam add_20099_20.INIT0 = 16'h5555;
    defparam add_20099_20.INIT1 = 16'h5555;
    defparam add_20099_20.INJECT1_0 = "NO";
    defparam add_20099_20.INJECT1_1 = "NO";
    CCU2D add_20099_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27503), .COUT(n27504));
    defparam add_20099_18.INIT0 = 16'h5555;
    defparam add_20099_18.INIT1 = 16'h5555;
    defparam add_20099_18.INJECT1_0 = "NO";
    defparam add_20099_18.INJECT1_1 = "NO";
    CCU2D add_20099_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27502), .COUT(n27503));
    defparam add_20099_16.INIT0 = 16'h5aaa;
    defparam add_20099_16.INIT1 = 16'h5555;
    defparam add_20099_16.INJECT1_0 = "NO";
    defparam add_20099_16.INJECT1_1 = "NO";
    CCU2D add_20099_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27501), .COUT(n27502));
    defparam add_20099_14.INIT0 = 16'h5aaa;
    defparam add_20099_14.INIT1 = 16'h5555;
    defparam add_20099_14.INJECT1_0 = "NO";
    defparam add_20099_14.INJECT1_1 = "NO";
    CCU2D add_20099_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27500), .COUT(n27501));
    defparam add_20099_12.INIT0 = 16'h5555;
    defparam add_20099_12.INIT1 = 16'h5aaa;
    defparam add_20099_12.INJECT1_0 = "NO";
    defparam add_20099_12.INJECT1_1 = "NO";
    CCU2D add_20099_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27499), .COUT(n27500));
    defparam add_20099_10.INIT0 = 16'h5aaa;
    defparam add_20099_10.INIT1 = 16'h5aaa;
    defparam add_20099_10.INJECT1_0 = "NO";
    defparam add_20099_10.INJECT1_1 = "NO";
    CCU2D add_20099_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27498), .COUT(n27499));
    defparam add_20099_8.INIT0 = 16'h5555;
    defparam add_20099_8.INIT1 = 16'h5aaa;
    defparam add_20099_8.INJECT1_0 = "NO";
    defparam add_20099_8.INJECT1_1 = "NO";
    CCU2D add_20099_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27497), .COUT(n27498));
    defparam add_20099_6.INIT0 = 16'h5555;
    defparam add_20099_6.INIT1 = 16'h5555;
    defparam add_20099_6.INJECT1_0 = "NO";
    defparam add_20099_6.INJECT1_1 = "NO";
    CCU2D add_20099_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27496), .COUT(n27497));
    defparam add_20099_4.INIT0 = 16'h5aaa;
    defparam add_20099_4.INIT1 = 16'h5aaa;
    defparam add_20099_4.INJECT1_0 = "NO";
    defparam add_20099_4.INJECT1_1 = "NO";
    CCU2D add_20099_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27496));
    defparam add_20099_2.INIT0 = 16'h7000;
    defparam add_20099_2.INIT1 = 16'h5555;
    defparam add_20099_2.INJECT1_0 = "NO";
    defparam add_20099_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module EncoderPeripheral_U11
//

module EncoderPeripheral_U11 (\read_size[0] , debug_c_c, n13797, n31923, 
            n27946, prev_select, n32001, read_value, \read_size[2] , 
            n15, \register_addr[0] , n31952, \quadA_delayed[2] , \quadB_delayed[1] , 
            n13779, encoder_li_c, encoder_lb_c, encoder_la_c, VCC_net, 
            GND_net, \quadA_delayed[1] , \quadB_delayed[2] ) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n13797;
    input n31923;
    input n27946;
    output prev_select;
    input n32001;
    output [31:0]read_value;
    output \read_size[2] ;
    input n15;
    input \register_addr[0] ;
    input n31952;
    input \quadA_delayed[2] ;
    input \quadB_delayed[1] ;
    output n13779;
    input encoder_li_c;
    input encoder_lb_c;
    input encoder_la_c;
    input VCC_net;
    input GND_net;
    input \quadA_delayed[1] ;
    input \quadB_delayed[2] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n29807;
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    wire [31:0]n100;
    
    wire n29819, n29817, n29809, n29811, n29810, n29812, n29813, 
        n29821, n29815, n6, n29808, n29818;
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n6_adj_535;
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n14851;
    wire [31:0]n180;
    
    wire n29820, n29816, n29814;
    
    FD1P3IX read_size__i1 (.D(n27946), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3AX prev_select_126 (.D(n32001), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam prev_select_126.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29807), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_size__i2 (.D(n15), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i14901_2_lut (.A(\register[1] [31]), .B(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14901_2_lut.init = 16'h8888;
    FD1P3AX read_value__i24 (.D(n29819), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29817), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i14902_2_lut (.A(\register[1] [30]), .B(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14902_2_lut.init = 16'h8888;
    LUT4 i14903_2_lut (.A(\register[1] [29]), .B(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14903_2_lut.init = 16'h8888;
    LUT4 i14904_2_lut (.A(\register[1] [28]), .B(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14904_2_lut.init = 16'h8888;
    LUT4 i14905_2_lut (.A(\register[1] [27]), .B(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14905_2_lut.init = 16'h8888;
    LUT4 i14906_2_lut (.A(\register[1] [26]), .B(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14906_2_lut.init = 16'h8888;
    LUT4 i14907_2_lut (.A(\register[1] [23]), .B(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14907_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [21]), 
         .Z(n29807)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_457 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [24]), 
         .Z(n29819)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_457.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_458 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [25]), 
         .Z(n29817)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_458.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_459 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [0]), 
         .Z(n29809)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_459.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_460 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [4]), 
         .Z(n29811)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_460.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_461 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [5]), 
         .Z(n29810)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_461.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_462 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [6]), 
         .Z(n29812)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_462.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_463 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [7]), 
         .Z(n29813)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_463.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_464 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [8]), 
         .Z(n29821)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_464.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_465 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [9]), 
         .Z(n29815)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_465.init = 16'h2020;
    LUT4 i1_4_lut (.A(n31952), .B(\quadA_delayed[2] ), .C(n6), .D(\quadB_delayed[1] ), 
         .Z(n13779)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(63[18:35])
    defparam i1_4_lut.init = 16'hebbe;
    LUT4 i14908_2_lut (.A(\register[1] [22]), .B(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14908_2_lut.init = 16'h8888;
    FD1P3AX read_value__i0 (.D(n29809), .SP(n13797), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_466 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [10]), 
         .Z(n29808)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_466.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_467 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [11]), 
         .Z(n29818)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_467.init = 16'h2020;
    LUT4 i14909_2_lut (.A(\register[1] [20]), .B(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14909_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_468 (.A(n31952), .B(quadA_delayed[2]), .C(n6_adj_535), 
         .D(quadB_delayed[2]), .Z(n14851)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(63[18:35])
    defparam i1_4_lut_adj_468.init = 16'hebbe;
    FD1P3IX read_value__i1 (.D(n180[1]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n180[2]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n180[3]), .SP(n13797), .CD(n31923), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29811), .SP(n13797), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29810), .SP(n13797), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29812), .SP(n13797), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 i14910_2_lut (.A(\register[1] [19]), .B(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14910_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_469 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [12]), 
         .Z(n29820)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_469.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_470 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [13]), 
         .Z(n29816)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_470.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_471 (.A(\register_addr[0] ), .B(n31923), .C(\register[1] [14]), 
         .Z(n29814)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam i1_2_lut_3_lut_adj_471.init = 16'h2020;
    LUT4 i14913_2_lut (.A(\register[1] [18]), .B(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14913_2_lut.init = 16'h8888;
    LUT4 i14914_2_lut (.A(\register[1] [17]), .B(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14914_2_lut.init = 16'h8888;
    FD1P3AX read_value__i7 (.D(n29813), .SP(n13797), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_li_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n180[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_lb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n180[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_la_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n180[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 i14915_2_lut (.A(\register[1] [16]), .B(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14915_2_lut.init = 16'h8888;
    LUT4 i14916_2_lut (.A(\register[1] [15]), .B(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14916_2_lut.init = 16'h8888;
    FD1P3AX read_value__i8 (.D(n29821), .SP(n13797), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29815), .SP(n13797), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29808), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29818), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29820), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29816), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29814), .SP(n13797), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=675, LSE_RLINE=685 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i14.GSR = "ENABLED";
    QuadratureDecoder_U6 q (.\register[1] ({\register[1] }), .debug_c_c(debug_c_c), 
            .n31952(n31952), .VCC_net(VCC_net), .GND_net(GND_net), .encoder_lb_c(encoder_lb_c), 
            .n14851(n14851), .encoder_la_c(encoder_la_c), .\quadA_delayed[1] (\quadA_delayed[1] ), 
            .\quadB_delayed[2] (\quadB_delayed[2] ), .n6(n6), .n6_adj_266(n6_adj_535), 
            .\quadB_delayed[2]_adj_267 (quadB_delayed[2]), .\quadA_delayed[2] (quadA_delayed[2])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(93[20] 97[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder_U6
//

module QuadratureDecoder_U6 (\register[1] , debug_c_c, n31952, VCC_net, 
            GND_net, encoder_lb_c, n14851, encoder_la_c, \quadA_delayed[1] , 
            \quadB_delayed[2] , n6, n6_adj_266, \quadB_delayed[2]_adj_267 , 
            \quadA_delayed[2] ) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[1] ;
    input debug_c_c;
    input n31952;
    input VCC_net;
    input GND_net;
    input encoder_lb_c;
    input n14851;
    input encoder_la_c;
    input \quadA_delayed[1] ;
    input \quadB_delayed[2] ;
    output n6;
    output n6_adj_266;
    output \quadB_delayed[2]_adj_267 ;
    output \quadA_delayed[2] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    wire [31:0]n100;
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [31:0]n4335;
    
    wire n27494, n27493, n27492, n27491, n27490, n27489, n27488, 
        n27487, n27486, n27485, n27484, n27483, n27482, n27481, 
        n27480, n27479;
    
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_lb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    FD1P3IX count__i0 (.D(n100[0]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_la_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    FD1P3IX count__i31 (.D(n4335[31]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4335[30]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n4335[1]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(\quadA_delayed[1] ), .B(\quadB_delayed[2] ), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    defparam i2_2_lut.init = 16'h6666;
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    LUT4 i2_2_lut_adj_456 (.A(quadA_delayed[1]), .B(quadB_delayed[1]), .Z(n6_adj_266)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    defparam i2_2_lut_adj_456.init = 16'h6666;
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(quadB_delayed[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(quadB_delayed[1]), .CK(debug_c_c), .Q(\quadB_delayed[2]_adj_267 )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n100[2]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n100[3]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n100[4]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n100[5]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n100[6]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n100[7]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n100[8]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n100[9]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n100[10]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n100[11]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n100[12]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n100[13]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n100[14]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n100[15]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n100[16]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n100[17]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n100[18]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n100[19]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n100[20]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n100[21]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n100[22]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n100[23]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n100[24]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n100[25]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n100[26]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n100[27]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n100[28]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n100[29]), .SP(n14851), .CD(n31952), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed[0]), .CK(debug_c_c), .Q(quadA_delayed[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(quadA_delayed[1]), .CK(debug_c_c), .Q(\quadA_delayed[2] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    CCU2D add_1667_33 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[30]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[31]), .D1(GND_net), .CIN(n27494), 
          .S0(n4335[30]), .S1(n4335[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_33.INIT0 = 16'h6969;
    defparam add_1667_33.INIT1 = 16'h6969;
    defparam add_1667_33.INJECT1_0 = "NO";
    defparam add_1667_33.INJECT1_1 = "NO";
    CCU2D add_1667_31 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[28]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[29]), .D1(GND_net), .CIN(n27493), 
          .COUT(n27494), .S0(n100[28]), .S1(n100[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_31.INIT0 = 16'h6969;
    defparam add_1667_31.INIT1 = 16'h6969;
    defparam add_1667_31.INJECT1_0 = "NO";
    defparam add_1667_31.INJECT1_1 = "NO";
    CCU2D add_1667_29 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[26]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[27]), .D1(GND_net), .CIN(n27492), 
          .COUT(n27493), .S0(n100[26]), .S1(n100[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_29.INIT0 = 16'h6969;
    defparam add_1667_29.INIT1 = 16'h6969;
    defparam add_1667_29.INJECT1_0 = "NO";
    defparam add_1667_29.INJECT1_1 = "NO";
    CCU2D add_1667_27 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[24]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[25]), .D1(GND_net), .CIN(n27491), 
          .COUT(n27492), .S0(n100[24]), .S1(n100[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_27.INIT0 = 16'h6969;
    defparam add_1667_27.INIT1 = 16'h6969;
    defparam add_1667_27.INJECT1_0 = "NO";
    defparam add_1667_27.INJECT1_1 = "NO";
    CCU2D add_1667_25 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[22]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[23]), .D1(GND_net), .CIN(n27490), 
          .COUT(n27491), .S0(n100[22]), .S1(n100[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_25.INIT0 = 16'h6969;
    defparam add_1667_25.INIT1 = 16'h6969;
    defparam add_1667_25.INJECT1_0 = "NO";
    defparam add_1667_25.INJECT1_1 = "NO";
    CCU2D add_1667_23 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[20]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[21]), .D1(GND_net), .CIN(n27489), 
          .COUT(n27490), .S0(n100[20]), .S1(n100[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_23.INIT0 = 16'h6969;
    defparam add_1667_23.INIT1 = 16'h6969;
    defparam add_1667_23.INJECT1_0 = "NO";
    defparam add_1667_23.INJECT1_1 = "NO";
    CCU2D add_1667_21 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[18]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[19]), .D1(GND_net), .CIN(n27488), 
          .COUT(n27489), .S0(n100[18]), .S1(n100[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_21.INIT0 = 16'h6969;
    defparam add_1667_21.INIT1 = 16'h6969;
    defparam add_1667_21.INJECT1_0 = "NO";
    defparam add_1667_21.INJECT1_1 = "NO";
    CCU2D add_1667_19 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[16]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[17]), .D1(GND_net), .CIN(n27487), 
          .COUT(n27488), .S0(n100[16]), .S1(n100[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_19.INIT0 = 16'h6969;
    defparam add_1667_19.INIT1 = 16'h6969;
    defparam add_1667_19.INJECT1_0 = "NO";
    defparam add_1667_19.INJECT1_1 = "NO";
    CCU2D add_1667_17 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[14]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[15]), .D1(GND_net), .CIN(n27486), 
          .COUT(n27487), .S0(n100[14]), .S1(n100[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_17.INIT0 = 16'h6969;
    defparam add_1667_17.INIT1 = 16'h6969;
    defparam add_1667_17.INJECT1_0 = "NO";
    defparam add_1667_17.INJECT1_1 = "NO";
    CCU2D add_1667_15 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[12]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[13]), .D1(GND_net), .CIN(n27485), 
          .COUT(n27486), .S0(n100[12]), .S1(n100[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_15.INIT0 = 16'h6969;
    defparam add_1667_15.INIT1 = 16'h6969;
    defparam add_1667_15.INJECT1_0 = "NO";
    defparam add_1667_15.INJECT1_1 = "NO";
    CCU2D add_1667_13 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[10]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[11]), .D1(GND_net), .CIN(n27484), 
          .COUT(n27485), .S0(n100[10]), .S1(n100[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_13.INIT0 = 16'h6969;
    defparam add_1667_13.INIT1 = 16'h6969;
    defparam add_1667_13.INJECT1_0 = "NO";
    defparam add_1667_13.INJECT1_1 = "NO";
    CCU2D add_1667_11 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[8]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[9]), .D1(GND_net), .CIN(n27483), 
          .COUT(n27484), .S0(n100[8]), .S1(n100[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_11.INIT0 = 16'h6969;
    defparam add_1667_11.INIT1 = 16'h6969;
    defparam add_1667_11.INJECT1_0 = "NO";
    defparam add_1667_11.INJECT1_1 = "NO";
    CCU2D add_1667_9 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[6]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[7]), .D1(GND_net), .CIN(n27482), 
          .COUT(n27483), .S0(n100[6]), .S1(n100[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_9.INIT0 = 16'h6969;
    defparam add_1667_9.INIT1 = 16'h6969;
    defparam add_1667_9.INJECT1_0 = "NO";
    defparam add_1667_9.INJECT1_1 = "NO";
    CCU2D add_1667_7 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[4]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[5]), .D1(GND_net), .CIN(n27481), 
          .COUT(n27482), .S0(n100[4]), .S1(n100[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_7.INIT0 = 16'h6969;
    defparam add_1667_7.INIT1 = 16'h6969;
    defparam add_1667_7.INJECT1_0 = "NO";
    defparam add_1667_7.INJECT1_1 = "NO";
    CCU2D add_1667_5 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[2]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[3]), .D1(GND_net), .CIN(n27480), 
          .COUT(n27481), .S0(n100[2]), .S1(n100[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_5.INIT0 = 16'h6969;
    defparam add_1667_5.INIT1 = 16'h6969;
    defparam add_1667_5.INJECT1_0 = "NO";
    defparam add_1667_5.INJECT1_1 = "NO";
    CCU2D add_1667_3 (.A0(\quadB_delayed[2]_adj_267 ), .B0(quadA_delayed[1]), 
          .C0(count[0]), .D0(GND_net), .A1(\quadB_delayed[2]_adj_267 ), 
          .B1(quadA_delayed[1]), .C1(count[1]), .D1(GND_net), .CIN(n27479), 
          .COUT(n27480), .S0(n100[0]), .S1(n4335[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_3.INIT0 = 16'h9696;
    defparam add_1667_3.INIT1 = 16'h6969;
    defparam add_1667_3.INJECT1_0 = "NO";
    defparam add_1667_3.INJECT1_1 = "NO";
    CCU2D add_1667_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\quadB_delayed[2]_adj_267 ), .B1(quadA_delayed[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27479));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1667_1.INIT0 = 16'hF000;
    defparam add_1667_1.INIT1 = 16'h6666;
    defparam add_1667_1.INJECT1_0 = "NO";
    defparam add_1667_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (databus_out, n33683, read_value, read_value_adj_264, 
            n52, n46, n3, databus, \read_value[16]_adj_83 , read_value_adj_265, 
            n31924, n47, \read_value[16]_adj_116 , n6, n31942, n3_adj_117, 
            \read_value[15]_adj_118 , \read_value[15]_adj_119 , n6_adj_120, 
            rw, \register_addr[0] , n3_adj_121, \read_value[14]_adj_122 , 
            \read_value[14]_adj_123 , n6_adj_124, \select[7] , n3_adj_125, 
            \read_value[13]_adj_126 , \read_value[13]_adj_127 , n6_adj_128, 
            n3_adj_129, \read_value[30]_adj_130 , \read_value[30]_adj_131 , 
            n6_adj_132, n3_adj_133, \read_value[12]_adj_134 , \read_value[12]_adj_135 , 
            n6_adj_136, n3_adj_137, \read_value[29]_adj_138 , \read_value[29]_adj_139 , 
            n6_adj_140, n3_adj_141, \read_value[28]_adj_142 , \read_value[28]_adj_143 , 
            n6_adj_144, n3_adj_145, \read_value[27]_adj_146 , \read_value[27]_adj_147 , 
            n6_adj_148, n3_adj_149, \read_value[11]_adj_150 , \read_value[11]_adj_151 , 
            n6_adj_152, \register_addr[2] , n3_adj_153, \read_value[26]_adj_154 , 
            \read_value[26]_adj_155 , n6_adj_156, n3_adj_157, \read_value[10]_adj_158 , 
            \read_value[10]_adj_159 , n6_adj_160, \read_value[0]_adj_161 , 
            n31944, n3_adj_162, \read_value[9]_adj_163 , \read_value[9]_adj_164 , 
            n6_adj_165, \read_value[0]_adj_166 , read_size, \select[1] , 
            n32068, \sendcount[1] , n12930, n3_adj_167, \read_value[8]_adj_168 , 
            n3_adj_169, \read_value[25]_adj_170 , \read_value[25]_adj_171 , 
            n6_adj_172, \read_value[8]_adj_173 , n6_adj_174, \read_value[7]_adj_175 , 
            n5, n8, n3_adj_176, \read_value[24]_adj_177 , \read_value[24]_adj_178 , 
            n6_adj_179, \register_addr[1] , \read_value[7]_adj_180 , \read_value[7]_adj_181 , 
            n3_adj_182, \read_value[23]_adj_183 , \read_value[23]_adj_184 , 
            n6_adj_185, n3_adj_186, \read_value[22]_adj_187 , \read_value[22]_adj_188 , 
            n6_adj_189, n3_adj_190, \read_value[21]_adj_191 , \read_value[21]_adj_192 , 
            n6_adj_193, n3_adj_194, \read_value[20]_adj_195 , \read_value[20]_adj_196 , 
            n6_adj_197, n3_adj_198, \read_value[19]_adj_199 , \read_value[19]_adj_200 , 
            n6_adj_201, n32090, \register_addr[3] , n32089, n31987, 
            n13323, n31970, \register_addr[5] , n31972, n33680, n31975, 
            n3_adj_202, n32034, n32006, \read_value[18]_adj_203 , \read_value[18]_adj_204 , 
            n6_adj_205, n31965, \select[4] , \read_size[0]_adj_206 , 
            n22, \read_size[0]_adj_207 , n8_adj_208, \select[2] , n12, 
            n31990, \read_size[0]_adj_209 , n8_adj_210, \read_size[0]_adj_211 , 
            n30166, \read_size[0]_adj_212 , n31977, \read_size[0]_adj_213 , 
            n3_adj_214, \read_value[17]_adj_215 , \read_value[17]_adj_216 , 
            n6_adj_217, \reg_size[2] , \read_size[2]_adj_218 , n32001, 
            \read_size[2]_adj_219 , \read_size[2]_adj_220 , \read_size[2]_adj_221 , 
            \read_size[2]_adj_222 , \read_size[2]_adj_223 , \read_value[6]_adj_224 , 
            n5_adj_225, n8_adj_226, \read_value[6]_adj_227 , n4, \read_value[6]_adj_228 , 
            \read_value[1]_adj_229 , n31959, \read_value[5]_adj_230 , 
            n5_adj_231, n8_adj_232, \read_value[5]_adj_233 , \read_value[5]_adj_234 , 
            n32004, \read_value[4]_adj_235 , n5_adj_236, n1, n5_adj_237, 
            n8_adj_238, \read_value[4]_adj_239 , \read_value[4]_adj_240 , 
            \read_value[3]_adj_241 , n5_adj_242, n8_adj_243, \read_value[3]_adj_244 , 
            \read_value[3]_adj_245 , \read_value[2]_adj_246 , n5_adj_247, 
            \read_value[1]_adj_248 , n3_adj_249, \read_value[31]_adj_250 , 
            \read_value[31]_adj_251 , n6_adj_252, n8_adj_253, \read_value[2]_adj_254 , 
            \read_value[0]_adj_255 , n5_adj_256, \read_value[2]_adj_257 , 
            n8_adj_258, n32039, n5_adj_259, n27979, GND_net, debug_c_c, 
            n33686, rc_ch8_c, n30381, n33685, n13735, n27956, n27877, 
            rc_ch7_c, n5_adj_260, n32074, n28044, n27887, n27759, 
            n33687, n14315, n30505, \count[8] , \count[13] , n27644, 
            rc_ch4_c, \count[11] , n30520, \count[9] , \count[10] , 
            n32025, n154, n27883, n29469, n30220, n5_adj_261, n27879, 
            n30196, n27809, \count[8]_adj_262 , n30202, \count[9]_adj_263 , 
            \count[6] , \count[7] , n32062, \count[5] , n27853, n32064, 
            n27983, rc_ch3_c, n32080, n27758, n29341, n14358, n30445, 
            n1168, n1180, n31964, n30426, n31906, n14369, n27757, 
            rc_ch2_c, n29866, n1153, n1165, n31948, n30378, n14374, 
            rc_ch1_c, n27960, n29869) /* synthesis syn_module_defined=1 */ ;
    input [31:0]databus_out;
    input n33683;
    input [31:0]read_value;
    input [31:0]read_value_adj_264;
    input n52;
    input n46;
    input n3;
    output [31:0]databus;
    input \read_value[16]_adj_83 ;
    input [31:0]read_value_adj_265;
    input n31924;
    input n47;
    input \read_value[16]_adj_116 ;
    input n6;
    input n31942;
    input n3_adj_117;
    input \read_value[15]_adj_118 ;
    input \read_value[15]_adj_119 ;
    input n6_adj_120;
    input rw;
    input \register_addr[0] ;
    input n3_adj_121;
    input \read_value[14]_adj_122 ;
    input \read_value[14]_adj_123 ;
    input n6_adj_124;
    input \select[7] ;
    input n3_adj_125;
    input \read_value[13]_adj_126 ;
    input \read_value[13]_adj_127 ;
    input n6_adj_128;
    input n3_adj_129;
    input \read_value[30]_adj_130 ;
    input \read_value[30]_adj_131 ;
    input n6_adj_132;
    input n3_adj_133;
    input \read_value[12]_adj_134 ;
    input \read_value[12]_adj_135 ;
    input n6_adj_136;
    input n3_adj_137;
    input \read_value[29]_adj_138 ;
    input \read_value[29]_adj_139 ;
    input n6_adj_140;
    input n3_adj_141;
    input \read_value[28]_adj_142 ;
    input \read_value[28]_adj_143 ;
    input n6_adj_144;
    input n3_adj_145;
    input \read_value[27]_adj_146 ;
    input \read_value[27]_adj_147 ;
    input n6_adj_148;
    input n3_adj_149;
    input \read_value[11]_adj_150 ;
    input \read_value[11]_adj_151 ;
    input n6_adj_152;
    input \register_addr[2] ;
    input n3_adj_153;
    input \read_value[26]_adj_154 ;
    input \read_value[26]_adj_155 ;
    input n6_adj_156;
    input n3_adj_157;
    input \read_value[10]_adj_158 ;
    input \read_value[10]_adj_159 ;
    input n6_adj_160;
    input \read_value[0]_adj_161 ;
    input n31944;
    input n3_adj_162;
    input \read_value[9]_adj_163 ;
    input \read_value[9]_adj_164 ;
    input n6_adj_165;
    input \read_value[0]_adj_166 ;
    input [2:0]read_size;
    input \select[1] ;
    output n32068;
    input \sendcount[1] ;
    output n12930;
    input n3_adj_167;
    input \read_value[8]_adj_168 ;
    input n3_adj_169;
    input \read_value[25]_adj_170 ;
    input \read_value[25]_adj_171 ;
    input n6_adj_172;
    input \read_value[8]_adj_173 ;
    input n6_adj_174;
    input \read_value[7]_adj_175 ;
    input n5;
    input n8;
    input n3_adj_176;
    input \read_value[24]_adj_177 ;
    input \read_value[24]_adj_178 ;
    input n6_adj_179;
    input \register_addr[1] ;
    input \read_value[7]_adj_180 ;
    input \read_value[7]_adj_181 ;
    input n3_adj_182;
    input \read_value[23]_adj_183 ;
    input \read_value[23]_adj_184 ;
    input n6_adj_185;
    input n3_adj_186;
    input \read_value[22]_adj_187 ;
    input \read_value[22]_adj_188 ;
    input n6_adj_189;
    input n3_adj_190;
    input \read_value[21]_adj_191 ;
    input \read_value[21]_adj_192 ;
    input n6_adj_193;
    input n3_adj_194;
    input \read_value[20]_adj_195 ;
    input \read_value[20]_adj_196 ;
    input n6_adj_197;
    input n3_adj_198;
    input \read_value[19]_adj_199 ;
    input \read_value[19]_adj_200 ;
    input n6_adj_201;
    input n32090;
    input \register_addr[3] ;
    input n32089;
    output n31987;
    input n13323;
    output n31970;
    input \register_addr[5] ;
    output n31972;
    input n33680;
    output n31975;
    input n3_adj_202;
    input n32034;
    output n32006;
    input \read_value[18]_adj_203 ;
    input \read_value[18]_adj_204 ;
    input n6_adj_205;
    output n31965;
    input \select[4] ;
    input \read_size[0]_adj_206 ;
    output n22;
    input \read_size[0]_adj_207 ;
    input n8_adj_208;
    input \select[2] ;
    output n12;
    input n31990;
    input \read_size[0]_adj_209 ;
    output n8_adj_210;
    input \read_size[0]_adj_211 ;
    input n30166;
    input \read_size[0]_adj_212 ;
    input n31977;
    input \read_size[0]_adj_213 ;
    input n3_adj_214;
    input \read_value[17]_adj_215 ;
    input \read_value[17]_adj_216 ;
    input n6_adj_217;
    output \reg_size[2] ;
    input \read_size[2]_adj_218 ;
    input n32001;
    input \read_size[2]_adj_219 ;
    input \read_size[2]_adj_220 ;
    input \read_size[2]_adj_221 ;
    input \read_size[2]_adj_222 ;
    input \read_size[2]_adj_223 ;
    input \read_value[6]_adj_224 ;
    input n5_adj_225;
    input n8_adj_226;
    input \read_value[6]_adj_227 ;
    input n4;
    input \read_value[6]_adj_228 ;
    input \read_value[1]_adj_229 ;
    input n31959;
    input \read_value[5]_adj_230 ;
    input n5_adj_231;
    input n8_adj_232;
    input \read_value[5]_adj_233 ;
    input \read_value[5]_adj_234 ;
    input n32004;
    input \read_value[4]_adj_235 ;
    input n5_adj_236;
    input n1;
    input n5_adj_237;
    input n8_adj_238;
    input \read_value[4]_adj_239 ;
    input \read_value[4]_adj_240 ;
    input \read_value[3]_adj_241 ;
    input n5_adj_242;
    input n8_adj_243;
    input \read_value[3]_adj_244 ;
    input \read_value[3]_adj_245 ;
    input \read_value[2]_adj_246 ;
    input n5_adj_247;
    input \read_value[1]_adj_248 ;
    input n3_adj_249;
    input \read_value[31]_adj_250 ;
    input \read_value[31]_adj_251 ;
    input n6_adj_252;
    input n8_adj_253;
    input \read_value[2]_adj_254 ;
    input \read_value[0]_adj_255 ;
    input n5_adj_256;
    input \read_value[2]_adj_257 ;
    input n8_adj_258;
    output n32039;
    output n5_adj_259;
    output n27979;
    input GND_net;
    input debug_c_c;
    input n33686;
    input rc_ch8_c;
    output n30381;
    input n33685;
    input n13735;
    input n27956;
    output n27877;
    input rc_ch7_c;
    output n5_adj_260;
    output n32074;
    output n28044;
    output n27887;
    input n27759;
    input n33687;
    input n14315;
    output n30505;
    output \count[8] ;
    output \count[13] ;
    output n27644;
    input rc_ch4_c;
    output \count[11] ;
    output n30520;
    output \count[9] ;
    output \count[10] ;
    output n32025;
    output n154;
    input n27883;
    input n29469;
    input n30220;
    output n5_adj_261;
    output n27879;
    output n30196;
    output n27809;
    output \count[8]_adj_262 ;
    input n30202;
    output \count[9]_adj_263 ;
    output \count[6] ;
    output \count[7] ;
    output n32062;
    output \count[5] ;
    output n27853;
    output n32064;
    output n27983;
    input rc_ch3_c;
    output n32080;
    input n27758;
    input n29341;
    input n14358;
    output n30445;
    output n1168;
    output n1180;
    output n31964;
    output n30426;
    input n31906;
    input n14369;
    input n27757;
    input rc_ch2_c;
    output n29866;
    output n1153;
    output n1165;
    output n31948;
    output n30378;
    input n14374;
    input rc_ch1_c;
    input n27960;
    output n29869;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(461[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n5_c, n12_c, n9, n14, n5_adj_167, n12_adj_170, n9_adj_173, 
        n14_adj_174, n5_adj_176, n12_adj_179;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31026, n9_adj_183, n14_adj_184, n5_adj_186, n12_adj_189;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31669;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(211[12:21])
    
    wire n176;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31666, n31667, n1219;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31670, n9_adj_193, n14_adj_194, n5_adj_196, n12_adj_199, 
        n9_adj_201, n14_adj_202, n5_adj_204, n12_adj_209, n31006, 
        n31752, n9_adj_211, n14_adj_212, n5_adj_214, n12_adj_219, 
        n9_adj_221, n14_adj_222, n5_adj_224, n12_adj_227, n9_adj_231, 
        n14_adj_232, n5_adj_234, n12_adj_237, n9_adj_241, n14_adj_242, 
        n5_adj_244, n12_adj_247, n31755, n9_adj_251, n14_adj_252, 
        n5_adj_254, n31753, n31756, n12_adj_259, n31030, n31027, 
        n31031, n9_adj_261, n14_adj_262, n5_adj_264, n12_adj_269, 
        n31821, n9_adj_271, n14_adj_272, n5_adj_274, n12_adj_277, 
        n31822, n14_adj_284, n31824, n1159, n31825, n31841, n31840, 
        n31843, n1174, n31844, n9_adj_285, n14_adj_286, n5_adj_288, 
        n12_adj_291;
    wire [7:0]read_value_adj_529;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(210[12:22])
    
    wire n46_adj_295, n12_adj_296, n9_adj_299, n14_adj_300, n5_adj_302, 
        n9_adj_304, n14_adj_305, n5_adj_307, n12_adj_310, n12_adj_313, 
        n17, n6_adj_317, n16, n2, n31007, n14_adj_320, n12_adj_323, 
        n9_adj_324, n14_adj_325, n5_adj_327, n12_adj_330, n31029, 
        n31028, n1234, n31528, n31527, n31525, n31524, n9_adj_339, 
        n14_adj_340, n5_adj_342, n12_adj_345, n9_adj_349, n14_adj_350, 
        n5_adj_352, n12_adj_355, n9_adj_359, n14_adj_360, n5_adj_362, 
        n12_adj_365, n31586, n9_adj_369, n14_adj_370, n5_adj_372, 
        n12_adj_375, n9_adj_379, n14_adj_380, n5_adj_382, n31585, 
        n31588, n12_adj_385, n1189, n31589, n9_adj_389, n14_adj_390, 
        n5_adj_392, n12_adj_395, n29911, n10, n31025, n9_adj_409, 
        n14_adj_410, n7, n6_adj_416, n20, n17_adj_421, n1204, n17_adj_424, 
        n6_adj_425, n16_adj_426, n2_adj_427, n14_adj_428, n12_adj_431, 
        n11, n16_adj_436, n31004, n31949, n31846, n31591, n31758, 
        n31009, n31672, n31530, n31845, n31842, n2_adj_440, n31826, 
        n31823, n31827, n17_adj_441, n6_adj_442, n16_adj_443, n2_adj_444, 
        n31757, n31754, n14_adj_447, n31671, n31668, n12_adj_450, 
        n31003, n31590, n31587, n17_adj_456, n6_adj_457, n16_adj_458, 
        n2_adj_459, n14_adj_461, n31008, n18, n14_adj_463, n12_adj_467, 
        n31529, n31526, n17_adj_473, n6_adj_474, n16_adj_475, n2_adj_476, 
        n14_adj_478, n12_adj_481, n17_adj_487, n6_adj_488, n16_adj_489, 
        n2_adj_490, n14_adj_492, n31005, n9_adj_496, n14_adj_497, 
        n5_adj_499, n12_adj_502, n12_adj_505, n17_adj_508, n6_adj_509, 
        n16_adj_510, n2_adj_511;
    
    LUT4 Select_4219_i5_2_lut (.A(databus_out[17]), .B(n33683), .Z(n5_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4219_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut (.A(read_value[17]), .B(read_value_adj_264[17]), .C(n52), 
         .D(n46), .Z(n12_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut.init = 16'heca0;
    LUT4 i7_4_lut (.A(n9), .B(n14), .C(n3), .D(n5_adj_167), .Z(databus[16])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(\read_value[16]_adj_83 ), .B(read_value_adj_265[16]), 
         .C(n31924), .D(n47), .Z(n9)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i6_4_lut (.A(\read_value[16]_adj_116 ), .B(n12_adj_170), .C(n6), 
         .D(n31942), .Z(n14)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 Select_4222_i5_2_lut (.A(databus_out[16]), .B(n33683), .Z(n5_adj_167)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4222_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_320 (.A(read_value[16]), .B(read_value_adj_264[16]), 
         .C(n52), .D(n46), .Z(n12_adj_170)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_320.init = 16'heca0;
    LUT4 i7_4_lut_adj_321 (.A(n9_adj_173), .B(n14_adj_174), .C(n3_adj_117), 
         .D(n5_adj_176), .Z(databus[15])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_321.init = 16'hfffe;
    LUT4 i1_4_lut_adj_322 (.A(\read_value[15]_adj_118 ), .B(read_value_adj_265[15]), 
         .C(n31924), .D(n47), .Z(n9_adj_173)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_322.init = 16'heca0;
    LUT4 i6_4_lut_adj_323 (.A(\read_value[15]_adj_119 ), .B(n12_adj_179), 
         .C(n6_adj_120), .D(n31942), .Z(n14_adj_174)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_323.init = 16'hfefc;
    LUT4 Select_4225_i5_2_lut (.A(databus_out[15]), .B(rw), .Z(n5_adj_176)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4225_i5_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_23398 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n31026)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23398.init = 16'he4e4;
    LUT4 i4_4_lut_adj_324 (.A(read_value[15]), .B(read_value_adj_264[15]), 
         .C(n52), .D(n46), .Z(n12_adj_179)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_324.init = 16'heca0;
    LUT4 i7_4_lut_adj_325 (.A(n9_adj_183), .B(n14_adj_184), .C(n3_adj_121), 
         .D(n5_adj_186), .Z(databus[14])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_325.init = 16'hfffe;
    LUT4 i1_4_lut_adj_326 (.A(\read_value[14]_adj_122 ), .B(read_value_adj_265[14]), 
         .C(n31924), .D(n47), .Z(n9_adj_183)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_326.init = 16'heca0;
    LUT4 i6_4_lut_adj_327 (.A(\read_value[14]_adj_123 ), .B(n12_adj_189), 
         .C(n6_adj_124), .D(n31942), .Z(n14_adj_184)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_327.init = 16'hfefc;
    LUT4 Select_4228_i5_2_lut (.A(databus_out[14]), .B(rw), .Z(n5_adj_186)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4228_i5_2_lut.init = 16'h2222;
    LUT4 n1219_bdd_3_lut_23566 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n31669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1219_bdd_3_lut_23566.init = 16'hcaca;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 i4_4_lut_adj_328 (.A(read_value[14]), .B(read_value_adj_264[14]), 
         .C(n52), .D(n46), .Z(n12_adj_189)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_328.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_23581 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n31666)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23581.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_23582 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n31667)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23582.init = 16'he4e4;
    LUT4 n1219_bdd_3_lut_24062 (.A(n1219), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n31670)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1219_bdd_3_lut_24062.init = 16'he2e2;
    LUT4 i7_4_lut_adj_329 (.A(n9_adj_193), .B(n14_adj_194), .C(n3_adj_125), 
         .D(n5_adj_196), .Z(databus[13])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_329.init = 16'hfffe;
    LUT4 i1_4_lut_adj_330 (.A(\read_value[13]_adj_126 ), .B(read_value_adj_265[13]), 
         .C(n31924), .D(n47), .Z(n9_adj_193)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_330.init = 16'heca0;
    LUT4 i6_4_lut_adj_331 (.A(\read_value[13]_adj_127 ), .B(n12_adj_199), 
         .C(n6_adj_128), .D(n31942), .Z(n14_adj_194)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_331.init = 16'hfefc;
    LUT4 i7_4_lut_adj_332 (.A(n9_adj_201), .B(n14_adj_202), .C(n3_adj_129), 
         .D(n5_adj_204), .Z(databus[30])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_332.init = 16'hfffe;
    LUT4 i1_4_lut_adj_333 (.A(\read_value[30]_adj_130 ), .B(read_value_adj_265[30]), 
         .C(n31924), .D(n47), .Z(n9_adj_201)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_333.init = 16'heca0;
    LUT4 Select_4231_i5_2_lut (.A(databus_out[13]), .B(rw), .Z(n5_adj_196)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4231_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_334 (.A(read_value[13]), .B(read_value_adj_264[13]), 
         .C(n52), .D(n46), .Z(n12_adj_199)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_334.init = 16'heca0;
    LUT4 i6_4_lut_adj_335 (.A(\read_value[30]_adj_131 ), .B(n12_adj_209), 
         .C(n6_adj_132), .D(n31942), .Z(n14_adj_202)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_335.init = 16'hfefc;
    LUT4 Select_4180_i5_2_lut (.A(databus_out[30]), .B(rw), .Z(n5_adj_204)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4180_i5_2_lut.init = 16'h2222;
    LUT4 \register_1[[5__bdd_3_lut_23652  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n31006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_23652 .init = 16'hcaca;
    LUT4 register_addr_1__bdd_2_lut_23626 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n31752)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23626.init = 16'h2222;
    LUT4 i7_4_lut_adj_336 (.A(n9_adj_211), .B(n14_adj_212), .C(n3_adj_133), 
         .D(n5_adj_214), .Z(databus[12])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_336.init = 16'hfffe;
    LUT4 i4_4_lut_adj_337 (.A(read_value[30]), .B(read_value_adj_264[30]), 
         .C(n52), .D(n46), .Z(n12_adj_209)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_337.init = 16'heca0;
    LUT4 i1_4_lut_adj_338 (.A(\read_value[12]_adj_134 ), .B(read_value_adj_265[12]), 
         .C(n31924), .D(n47), .Z(n9_adj_211)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_338.init = 16'heca0;
    LUT4 i6_4_lut_adj_339 (.A(\read_value[12]_adj_135 ), .B(n12_adj_219), 
         .C(n6_adj_136), .D(n31942), .Z(n14_adj_212)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_339.init = 16'hfefc;
    LUT4 i7_4_lut_adj_340 (.A(n9_adj_221), .B(n14_adj_222), .C(n3_adj_137), 
         .D(n5_adj_224), .Z(databus[29])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_340.init = 16'hfffe;
    LUT4 i1_4_lut_adj_341 (.A(\read_value[29]_adj_138 ), .B(read_value_adj_265[29]), 
         .C(n31924), .D(n47), .Z(n9_adj_221)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_341.init = 16'heca0;
    LUT4 i6_4_lut_adj_342 (.A(\read_value[29]_adj_139 ), .B(n12_adj_227), 
         .C(n6_adj_140), .D(n31942), .Z(n14_adj_222)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_342.init = 16'hfefc;
    LUT4 Select_4183_i5_2_lut (.A(databus_out[29]), .B(rw), .Z(n5_adj_224)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4183_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_343 (.A(read_value[29]), .B(read_value_adj_264[29]), 
         .C(n52), .D(n46), .Z(n12_adj_227)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_343.init = 16'heca0;
    LUT4 i7_4_lut_adj_344 (.A(n9_adj_231), .B(n14_adj_232), .C(n3_adj_141), 
         .D(n5_adj_234), .Z(databus[28])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_344.init = 16'hfffe;
    LUT4 i1_4_lut_adj_345 (.A(\read_value[28]_adj_142 ), .B(read_value_adj_265[28]), 
         .C(n31924), .D(n47), .Z(n9_adj_231)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_345.init = 16'heca0;
    LUT4 i6_4_lut_adj_346 (.A(\read_value[28]_adj_143 ), .B(n12_adj_237), 
         .C(n6_adj_144), .D(n31942), .Z(n14_adj_232)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_346.init = 16'hfefc;
    LUT4 Select_4186_i5_2_lut (.A(databus_out[28]), .B(rw), .Z(n5_adj_234)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4186_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_347 (.A(read_value[28]), .B(read_value_adj_264[28]), 
         .C(n52), .D(n46), .Z(n12_adj_237)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_347.init = 16'heca0;
    LUT4 i7_4_lut_adj_348 (.A(n9_adj_241), .B(n14_adj_242), .C(n3_adj_145), 
         .D(n5_adj_244), .Z(databus[27])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_348.init = 16'hfffe;
    LUT4 i1_4_lut_adj_349 (.A(\read_value[27]_adj_146 ), .B(read_value_adj_265[27]), 
         .C(n31924), .D(n47), .Z(n9_adj_241)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_349.init = 16'heca0;
    LUT4 i6_4_lut_adj_350 (.A(\read_value[27]_adj_147 ), .B(n12_adj_247), 
         .C(n6_adj_148), .D(n31942), .Z(n14_adj_242)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_350.init = 16'hfefc;
    LUT4 Select_4234_i5_2_lut (.A(databus_out[12]), .B(rw), .Z(n5_adj_214)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4234_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_351 (.A(read_value[12]), .B(read_value_adj_264[12]), 
         .C(n52), .D(n46), .Z(n12_adj_219)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_351.init = 16'heca0;
    LUT4 \register_1[[4__bdd_3_lut_24010  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n31755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_24010 .init = 16'hcaca;
    LUT4 i7_4_lut_adj_352 (.A(n9_adj_251), .B(n14_adj_252), .C(n3_adj_149), 
         .D(n5_adj_254), .Z(databus[11])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_352.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_23627 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n31753)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23627.init = 16'he4e4;
    LUT4 i1_4_lut_adj_353 (.A(\read_value[11]_adj_150 ), .B(read_value_adj_265[11]), 
         .C(n31924), .D(n47), .Z(n9_adj_251)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_353.init = 16'heca0;
    LUT4 Select_4189_i5_2_lut (.A(databus_out[27]), .B(rw), .Z(n5_adj_244)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4189_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_354 (.A(read_value[27]), .B(read_value_adj_264[27]), 
         .C(n52), .D(n46), .Z(n12_adj_247)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_354.init = 16'heca0;
    LUT4 \register_1[[4__bdd_2_lut_24011  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n31756)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_24011 .init = 16'h8888;
    LUT4 i6_4_lut_adj_355 (.A(\read_value[11]_adj_151 ), .B(n12_adj_259), 
         .C(n6_adj_152), .D(n31942), .Z(n14_adj_252)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_355.init = 16'hfefc;
    L6MUX21 i23322 (.D0(n31030), .D1(n31027), .SD(\register_addr[2] ), 
            .Z(n31031));
    LUT4 i7_4_lut_adj_356 (.A(n9_adj_261), .B(n14_adj_262), .C(n3_adj_153), 
         .D(n5_adj_264), .Z(databus[26])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_356.init = 16'hfffe;
    LUT4 Select_4237_i5_2_lut (.A(databus_out[11]), .B(rw), .Z(n5_adj_254)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4237_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_357 (.A(read_value[11]), .B(read_value_adj_264[11]), 
         .C(n52), .D(n46), .Z(n12_adj_259)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_357.init = 16'heca0;
    LUT4 i1_4_lut_adj_358 (.A(\read_value[26]_adj_154 ), .B(read_value_adj_265[26]), 
         .C(n31924), .D(n47), .Z(n9_adj_261)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_358.init = 16'heca0;
    LUT4 i6_4_lut_adj_359 (.A(\read_value[26]_adj_155 ), .B(n12_adj_269), 
         .C(n6_adj_156), .D(n31942), .Z(n14_adj_262)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_359.init = 16'hfefc;
    LUT4 Select_4192_i5_2_lut (.A(databus_out[26]), .B(rw), .Z(n5_adj_264)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4192_i5_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_2_lut_23638 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n31821)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23638.init = 16'h2222;
    LUT4 i7_4_lut_adj_360 (.A(n9_adj_271), .B(n14_adj_272), .C(n3_adj_157), 
         .D(n5_adj_274), .Z(databus[10])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_360.init = 16'hfffe;
    LUT4 i1_4_lut_adj_361 (.A(\read_value[10]_adj_158 ), .B(read_value_adj_265[10]), 
         .C(n31924), .D(n47), .Z(n9_adj_271)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_361.init = 16'heca0;
    LUT4 i6_4_lut_adj_362 (.A(\read_value[10]_adj_159 ), .B(n12_adj_277), 
         .C(n6_adj_160), .D(n31942), .Z(n14_adj_272)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_362.init = 16'hfefc;
    LUT4 i4_4_lut_adj_363 (.A(read_value[26]), .B(read_value_adj_264[26]), 
         .C(n52), .D(n46), .Z(n12_adj_269)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_363.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23639 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n31822)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23639.init = 16'he4e4;
    LUT4 Select_4240_i5_2_lut (.A(databus_out[10]), .B(n33683), .Z(n5_adj_274)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4240_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_364 (.A(read_value[10]), .B(read_value_adj_264[10]), 
         .C(n52), .D(n46), .Z(n12_adj_277)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_364.init = 16'heca0;
    LUT4 i4_4_lut_adj_365 (.A(read_value_adj_264[0]), .B(\read_value[0]_adj_161 ), 
         .C(n46), .D(n31944), .Z(n14_adj_284)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_365.init = 16'heca0;
    LUT4 n1159_bdd_3_lut_23632 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n31824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1159_bdd_3_lut_23632.init = 16'hcaca;
    LUT4 n1159_bdd_3_lut_23929 (.A(n1159), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n31825)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1159_bdd_3_lut_23929.init = 16'he2e2;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n31841)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n31840)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    LUT4 n1174_bdd_3_lut_23645 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n31843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1174_bdd_3_lut_23645.init = 16'hcaca;
    LUT4 n1174_bdd_3_lut_23879 (.A(n1174), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n31844)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1174_bdd_3_lut_23879.init = 16'he2e2;
    LUT4 i7_4_lut_adj_366 (.A(n9_adj_285), .B(n14_adj_286), .C(n3_adj_162), 
         .D(n5_adj_288), .Z(databus[9])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_366.init = 16'hfffe;
    LUT4 i1_4_lut_adj_367 (.A(\read_value[9]_adj_163 ), .B(read_value_adj_265[9]), 
         .C(n31924), .D(n47), .Z(n9_adj_285)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_367.init = 16'heca0;
    LUT4 i6_4_lut_adj_368 (.A(\read_value[9]_adj_164 ), .B(n12_adj_291), 
         .C(n6_adj_165), .D(n31942), .Z(n14_adj_286)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_368.init = 16'hfefc;
    LUT4 i2_4_lut (.A(\read_value[0]_adj_166 ), .B(read_value_adj_529[0]), 
         .C(n31942), .D(n46_adj_295), .Z(n12_adj_296)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 Select_4243_i5_2_lut (.A(databus_out[9]), .B(rw), .Z(n5_adj_288)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4243_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_369 (.A(read_value[9]), .B(read_value_adj_264[9]), 
         .C(n52), .D(n46), .Z(n12_adj_291)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_369.init = 16'heca0;
    LUT4 Select_4263_i1_2_lut_rep_451 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n32068)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4263_i1_2_lut_rep_451.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n12930)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 i14_2_lut (.A(\select[7] ), .B(rw), .Z(n46_adj_295)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam i14_2_lut.init = 16'h8888;
    LUT4 i7_4_lut_adj_370 (.A(n9_adj_299), .B(n14_adj_300), .C(n3_adj_167), 
         .D(n5_adj_302), .Z(databus[8])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_370.init = 16'hfffe;
    LUT4 i1_4_lut_adj_371 (.A(\read_value[8]_adj_168 ), .B(read_value_adj_265[8]), 
         .C(n31924), .D(n47), .Z(n9_adj_299)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_371.init = 16'heca0;
    LUT4 i7_4_lut_adj_372 (.A(n9_adj_304), .B(n14_adj_305), .C(n3_adj_169), 
         .D(n5_adj_307), .Z(databus[25])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_372.init = 16'hfffe;
    LUT4 i1_4_lut_adj_373 (.A(\read_value[25]_adj_170 ), .B(read_value_adj_265[25]), 
         .C(n31924), .D(n47), .Z(n9_adj_304)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_373.init = 16'heca0;
    LUT4 i6_4_lut_adj_374 (.A(\read_value[25]_adj_171 ), .B(n12_adj_310), 
         .C(n6_adj_172), .D(n31942), .Z(n14_adj_305)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_374.init = 16'hfefc;
    LUT4 i6_4_lut_adj_375 (.A(\read_value[8]_adj_173 ), .B(n12_adj_313), 
         .C(n6_adj_174), .D(n31942), .Z(n14_adj_300)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_375.init = 16'hfefc;
    LUT4 Select_4195_i5_2_lut (.A(databus_out[25]), .B(rw), .Z(n5_adj_307)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4195_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_376 (.A(read_value[25]), .B(read_value_adj_264[25]), 
         .C(n52), .D(n46), .Z(n12_adj_310)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_376.init = 16'heca0;
    LUT4 i9_4_lut (.A(n17), .B(n6_adj_317), .C(n16), .D(n2), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 Select_4246_i5_2_lut (.A(databus_out[8]), .B(rw), .Z(n5_adj_302)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4246_i5_2_lut.init = 16'h2222;
    LUT4 \register_1[[5__bdd_2_lut_23653  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n31007)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_23653 .init = 16'h8888;
    LUT4 i4_4_lut_adj_377 (.A(read_value[8]), .B(read_value_adj_264[8]), 
         .C(n52), .D(n46), .Z(n12_adj_313)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_377.init = 16'heca0;
    LUT4 i7_4_lut_adj_378 (.A(\read_value[7]_adj_175 ), .B(n14_adj_320), 
         .C(n5), .D(n31924), .Z(n17)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_378.init = 16'hfefc;
    LUT4 Select_4247_i6_2_lut (.A(databus_out[7]), .B(rw), .Z(n6_adj_317)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4247_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_379 (.A(read_value_adj_265[7]), .B(n12_adj_323), .C(n8), 
         .D(n47), .Z(n16)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_379.init = 16'hfefc;
    LUT4 i7_4_lut_adj_380 (.A(n9_adj_324), .B(n14_adj_325), .C(n3_adj_176), 
         .D(n5_adj_327), .Z(databus[24])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_380.init = 16'hfffe;
    LUT4 i1_4_lut_adj_381 (.A(\read_value[24]_adj_177 ), .B(read_value_adj_265[24]), 
         .C(n31924), .D(n47), .Z(n9_adj_324)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_381.init = 16'heca0;
    LUT4 i6_4_lut_adj_382 (.A(\read_value[24]_adj_178 ), .B(n12_adj_330), 
         .C(n6_adj_179), .D(n31942), .Z(n14_adj_325)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_382.init = 16'hfefc;
    LUT4 Select_4198_i5_2_lut (.A(databus_out[24]), .B(rw), .Z(n5_adj_327)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4198_i5_2_lut.init = 16'h2222;
    LUT4 Select_4247_i2_2_lut (.A(read_value[7]), .B(n52), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4247_i2_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_383 (.A(read_value[24]), .B(read_value_adj_264[24]), 
         .C(n52), .D(n46), .Z(n12_adj_330)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_383.init = 16'heca0;
    PFUMX i23320 (.BLUT(n31029), .ALUT(n31028), .C0(\register_addr[1] ), 
          .Z(n31030));
    LUT4 i4_4_lut_adj_384 (.A(read_value_adj_264[7]), .B(\read_value[7]_adj_180 ), 
         .C(n46), .D(n31944), .Z(n14_adj_320)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_384.init = 16'heca0;
    LUT4 n1234_bdd_3_lut_23606 (.A(n1234), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n31528)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1234_bdd_3_lut_23606.init = 16'he2e2;
    LUT4 i2_4_lut_adj_385 (.A(\read_value[7]_adj_181 ), .B(read_value_adj_529[7]), 
         .C(n31942), .D(n46_adj_295), .Z(n12_adj_323)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_385.init = 16'heca0;
    LUT4 n1234_bdd_3_lut_23493 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n31527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1234_bdd_3_lut_23493.init = 16'hcaca;
    LUT4 register_addr_1__bdd_3_lut_23513 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n31525)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23513.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_23512 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n31524)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23512.init = 16'h2222;
    LUT4 i7_4_lut_adj_386 (.A(n9_adj_339), .B(n14_adj_340), .C(n3_adj_182), 
         .D(n5_adj_342), .Z(databus[23])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_386.init = 16'hfffe;
    LUT4 i1_4_lut_adj_387 (.A(\read_value[23]_adj_183 ), .B(read_value_adj_265[23]), 
         .C(n31924), .D(n47), .Z(n9_adj_339)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_387.init = 16'heca0;
    LUT4 i6_4_lut_adj_388 (.A(\read_value[23]_adj_184 ), .B(n12_adj_345), 
         .C(n6_adj_185), .D(n31942), .Z(n14_adj_340)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_388.init = 16'hfefc;
    LUT4 Select_4201_i5_2_lut (.A(databus_out[23]), .B(n33683), .Z(n5_adj_342)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4201_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_389 (.A(read_value[23]), .B(read_value_adj_264[23]), 
         .C(n52), .D(n46), .Z(n12_adj_345)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_389.init = 16'heca0;
    LUT4 i7_4_lut_adj_390 (.A(n9_adj_349), .B(n14_adj_350), .C(n3_adj_186), 
         .D(n5_adj_352), .Z(databus[22])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_390.init = 16'hfffe;
    LUT4 i1_4_lut_adj_391 (.A(\read_value[22]_adj_187 ), .B(read_value_adj_265[22]), 
         .C(n31924), .D(n47), .Z(n9_adj_349)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_391.init = 16'heca0;
    LUT4 i6_4_lut_adj_392 (.A(\read_value[22]_adj_188 ), .B(n12_adj_355), 
         .C(n6_adj_189), .D(n31942), .Z(n14_adj_350)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_392.init = 16'hfefc;
    LUT4 Select_4204_i5_2_lut (.A(databus_out[22]), .B(n33683), .Z(n5_adj_352)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4204_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_393 (.A(read_value[22]), .B(read_value_adj_264[22]), 
         .C(n52), .D(n46), .Z(n12_adj_355)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_393.init = 16'heca0;
    LUT4 i7_4_lut_adj_394 (.A(n9_adj_359), .B(n14_adj_360), .C(n3_adj_190), 
         .D(n5_adj_362), .Z(databus[21])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_394.init = 16'hfffe;
    LUT4 i1_4_lut_adj_395 (.A(\read_value[21]_adj_191 ), .B(read_value_adj_265[21]), 
         .C(n31924), .D(n47), .Z(n9_adj_359)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_395.init = 16'heca0;
    LUT4 i6_4_lut_adj_396 (.A(\read_value[21]_adj_192 ), .B(n12_adj_365), 
         .C(n6_adj_193), .D(n31942), .Z(n14_adj_360)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_396.init = 16'hfefc;
    LUT4 Select_4207_i5_2_lut (.A(databus_out[21]), .B(n33683), .Z(n5_adj_362)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4207_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_397 (.A(read_value[21]), .B(read_value_adj_264[21]), 
         .C(n52), .D(n46), .Z(n12_adj_365)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_397.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23561 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n31586)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23561.init = 16'he4e4;
    LUT4 i7_4_lut_adj_398 (.A(n9_adj_369), .B(n14_adj_370), .C(n3_adj_194), 
         .D(n5_adj_372), .Z(databus[20])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_398.init = 16'hfffe;
    LUT4 i1_4_lut_adj_399 (.A(\read_value[20]_adj_195 ), .B(read_value_adj_265[20]), 
         .C(n31924), .D(n47), .Z(n9_adj_369)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_399.init = 16'heca0;
    LUT4 i6_4_lut_adj_400 (.A(\read_value[20]_adj_196 ), .B(n12_adj_375), 
         .C(n6_adj_197), .D(n31942), .Z(n14_adj_370)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_400.init = 16'hfefc;
    LUT4 Select_4210_i5_2_lut (.A(databus_out[20]), .B(n33683), .Z(n5_adj_372)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4210_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_401 (.A(read_value[20]), .B(read_value_adj_264[20]), 
         .C(n52), .D(n46), .Z(n12_adj_375)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_401.init = 16'heca0;
    LUT4 i7_4_lut_adj_402 (.A(n9_adj_379), .B(n14_adj_380), .C(n3_adj_198), 
         .D(n5_adj_382), .Z(databus[19])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_402.init = 16'hfffe;
    LUT4 i1_4_lut_adj_403 (.A(\read_value[19]_adj_199 ), .B(read_value_adj_265[19]), 
         .C(n31924), .D(n47), .Z(n9_adj_379)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_403.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_23560 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n31585)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23560.init = 16'h2222;
    LUT4 n1189_bdd_3_lut_23524 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n31588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1189_bdd_3_lut_23524.init = 16'hcaca;
    LUT4 i6_4_lut_adj_404 (.A(\read_value[19]_adj_200 ), .B(n12_adj_385), 
         .C(n6_adj_201), .D(n31942), .Z(n14_adj_380)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_404.init = 16'hfefc;
    LUT4 i1_3_lut_rep_370_4_lut (.A(n32090), .B(\register_addr[3] ), .C(n32089), 
         .D(\register_addr[1] ), .Z(n31987)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_3_lut_rep_370_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_353_3_lut_4_lut (.A(n32090), .B(\register_addr[3] ), 
         .C(n13323), .D(\register_addr[2] ), .Z(n31970)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_353_3_lut_4_lut.init = 16'h0010;
    LUT4 n1189_bdd_3_lut_23573 (.A(n1189), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n31589)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1189_bdd_3_lut_23573.init = 16'he2e2;
    LUT4 Select_4213_i5_2_lut (.A(databus_out[19]), .B(n33683), .Z(n5_adj_382)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4213_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_405 (.A(read_value[19]), .B(read_value_adj_264[19]), 
         .C(n52), .D(n46), .Z(n12_adj_385)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_405.init = 16'heca0;
    LUT4 i1_2_lut_rep_355_3_lut_4_lut (.A(n32090), .B(\register_addr[3] ), 
         .C(\register_addr[5] ), .D(\register_addr[2] ), .Z(n31972)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_355_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_358_3_lut_4_lut (.A(n32090), .B(\register_addr[3] ), 
         .C(n33680), .D(\register_addr[2] ), .Z(n31975)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_358_3_lut_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut_adj_406 (.A(n9_adj_389), .B(n14_adj_390), .C(n3_adj_202), 
         .D(n5_adj_392), .Z(databus[18])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_406.init = 16'hfffe;
    LUT4 i22760_3_lut_rep_389_4_lut (.A(n32090), .B(\register_addr[3] ), 
         .C(\register_addr[5] ), .D(n32034), .Z(n32006)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22760_3_lut_rep_389_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_407 (.A(\read_value[18]_adj_203 ), .B(read_value_adj_265[18]), 
         .C(n31924), .D(n47), .Z(n9_adj_389)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_407.init = 16'heca0;
    LUT4 i6_4_lut_adj_408 (.A(\read_value[18]_adj_204 ), .B(n12_adj_395), 
         .C(n6_adj_205), .D(n31942), .Z(n14_adj_390)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_408.init = 16'hfefc;
    LUT4 i1_2_lut_rep_348_3_lut_4_lut (.A(n32090), .B(\register_addr[3] ), 
         .C(\register_addr[2] ), .D(n33680), .Z(n31965)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_348_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_409 (.A(\select[4] ), .B(\read_size[0]_adj_206 ), 
         .C(n29911), .D(n31970), .Z(n22)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_409.init = 16'ha8a0;
    LUT4 i5_4_lut (.A(\read_size[0]_adj_207 ), .B(n10), .C(n8_adj_208), 
         .D(\select[2] ), .Z(n12)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfefc;
    LUT4 i1_4_lut_adj_410 (.A(n31990), .B(\select[7] ), .C(\read_size[0]_adj_209 ), 
         .D(read_size_c[0]), .Z(n8_adj_210)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_410.init = 16'heca0;
    LUT4 Select_4216_i5_2_lut (.A(databus_out[18]), .B(n33683), .Z(n5_adj_392)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4216_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_411 (.A(read_value[18]), .B(read_value_adj_264[18]), 
         .C(n52), .D(n46), .Z(n12_adj_395)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_411.init = 16'heca0;
    LUT4 i1_4_lut_adj_412 (.A(\read_size[0]_adj_211 ), .B(n30166), .C(\read_size[0]_adj_212 ), 
         .D(\register_addr[5] ), .Z(n29911)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_412.init = 16'h3022;
    LUT4 i3_4_lut (.A(read_size[0]), .B(n31977), .C(\select[1] ), .D(\read_size[0]_adj_213 ), 
         .Z(n10)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_23397 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n31025)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23397.init = 16'h2222;
    LUT4 i7_4_lut_adj_413 (.A(n9_adj_409), .B(n14_adj_410), .C(n3_adj_214), 
         .D(n5_c), .Z(databus[17])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_413.init = 16'hfffe;
    LUT4 i1_4_lut_adj_414 (.A(\read_value[17]_adj_215 ), .B(read_value_adj_265[17]), 
         .C(n31924), .D(n47), .Z(n9_adj_409)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_414.init = 16'heca0;
    LUT4 i6_4_lut_adj_415 (.A(\read_value[17]_adj_216 ), .B(n12_c), .C(n6_adj_217), 
         .D(n31942), .Z(n14_adj_410)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_415.init = 16'hfefc;
    LUT4 i4_4_lut_adj_416 (.A(n7), .B(\select[4] ), .C(n6_adj_416), .D(n20), 
         .Z(\reg_size[2] )) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_416.init = 16'hfefa;
    LUT4 n1204_bdd_3_lut_23319 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n31028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1204_bdd_3_lut_23319.init = 16'hcaca;
    LUT4 i2_4_lut_adj_417 (.A(\read_size[2]_adj_218 ), .B(n31977), .C(n32001), 
         .D(\read_size[2]_adj_219 ), .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_417.init = 16'heca0;
    LUT4 i1_4_lut_adj_418 (.A(\select[1] ), .B(\read_size[2]_adj_220 ), 
         .C(read_size[2]), .D(n31990), .Z(n6_adj_416)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_418.init = 16'heca0;
    LUT4 i1_4_lut_adj_419 (.A(\read_size[2]_adj_221 ), .B(n17_adj_421), 
         .C(n31970), .D(n30166), .Z(n20)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam i1_4_lut_adj_419.init = 16'ha0ec;
    LUT4 i31_3_lut (.A(\read_size[2]_adj_222 ), .B(\read_size[2]_adj_223 ), 
         .C(\register_addr[5] ), .Z(n17_adj_421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31_3_lut.init = 16'hcaca;
    LUT4 n1204_bdd_3_lut_23326 (.A(n1204), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n31029)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1204_bdd_3_lut_23326.init = 16'he2e2;
    LUT4 i9_4_lut_adj_420 (.A(n17_adj_424), .B(n6_adj_425), .C(n16_adj_426), 
         .D(n2_adj_427), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_420.init = 16'hfffe;
    LUT4 i7_4_lut_adj_421 (.A(\read_value[6]_adj_224 ), .B(n14_adj_428), 
         .C(n5_adj_225), .D(n31924), .Z(n17_adj_424)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_421.init = 16'hfefc;
    LUT4 Select_4248_i6_2_lut (.A(databus_out[6]), .B(rw), .Z(n6_adj_425)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4248_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_422 (.A(read_value_adj_265[6]), .B(n12_adj_431), .C(n8_adj_226), 
         .D(n47), .Z(n16_adj_426)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_422.init = 16'hfefc;
    LUT4 Select_4248_i2_2_lut (.A(read_value[6]), .B(n52), .Z(n2_adj_427)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4248_i2_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_423 (.A(read_value_adj_264[6]), .B(\read_value[6]_adj_227 ), 
         .C(n46), .D(n31944), .Z(n14_adj_428)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_423.init = 16'heca0;
    LUT4 i6_4_lut_adj_424 (.A(n11), .B(n4), .C(databus_out[1]), .D(rw), 
         .Z(n16_adj_436)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i6_4_lut_adj_424.init = 16'heefe;
    LUT4 register_addr_1__bdd_3_lut_23316 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n31004)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23316.init = 16'he4e4;
    FD1S3IX read_value__i1 (.D(n31846), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n31591), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n31031), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n31758), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n31009), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(n31672), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i7 (.D(n31530), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_425 (.A(\read_value[6]_adj_228 ), .B(read_value_adj_529[6]), 
         .C(n31942), .D(n46_adj_295), .Z(n12_adj_431)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_425.init = 16'heca0;
    L6MUX21 i23648 (.D0(n31845), .D1(n31842), .SD(\register_addr[2] ), 
            .Z(n31846));
    PFUMX i23646 (.BLUT(n31844), .ALUT(n31843), .C0(\register_addr[1] ), 
          .Z(n31845));
    LUT4 Select_4253_i2_2_lut (.A(read_value[1]), .B(n52), .Z(n2_adj_440)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4253_i2_2_lut.init = 16'h8888;
    PFUMX i23643 (.BLUT(n31841), .ALUT(n31840), .C0(\register_addr[1] ), 
          .Z(n31842));
    L6MUX21 i23635 (.D0(n31826), .D1(n31823), .SD(\register_addr[2] ), 
            .Z(n31827));
    PFUMX i23633 (.BLUT(n31825), .ALUT(n31824), .C0(\register_addr[1] ), 
          .Z(n31826));
    PFUMX i23630 (.BLUT(n31822), .ALUT(n31821), .C0(\register_addr[1] ), 
          .Z(n31823));
    LUT4 i9_4_lut_adj_426 (.A(n17_adj_441), .B(n6_adj_442), .C(n16_adj_443), 
         .D(n2_adj_444), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_426.init = 16'hfffe;
    LUT4 i1_4_lut_adj_427 (.A(\read_value[1]_adj_229 ), .B(read_value_adj_529[1]), 
         .C(n31959), .D(n46_adj_295), .Z(n11)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_427.init = 16'heca0;
    L6MUX21 i23589 (.D0(n31757), .D1(n31754), .SD(\register_addr[2] ), 
            .Z(n31758));
    PFUMX i23587 (.BLUT(n31756), .ALUT(n31755), .C0(\register_addr[1] ), 
          .Z(n31757));
    PFUMX i23317 (.BLUT(n31026), .ALUT(n31025), .C0(\register_addr[1] ), 
          .Z(n31027));
    PFUMX i23585 (.BLUT(n31753), .ALUT(n31752), .C0(\register_addr[1] ), 
          .Z(n31754));
    LUT4 i7_4_lut_adj_428 (.A(\read_value[5]_adj_230 ), .B(n14_adj_447), 
         .C(n5_adj_231), .D(n31924), .Z(n17_adj_441)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_428.init = 16'hfefc;
    LUT4 Select_4249_i6_2_lut (.A(databus_out[5]), .B(n33683), .Z(n6_adj_442)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4249_i6_2_lut.init = 16'h2222;
    L6MUX21 i23569 (.D0(n31671), .D1(n31668), .SD(\register_addr[2] ), 
            .Z(n31672));
    LUT4 i6_4_lut_adj_429 (.A(read_value_adj_265[5]), .B(n12_adj_450), .C(n8_adj_232), 
         .D(n47), .Z(n16_adj_443)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_429.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_23315 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n31003)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23315.init = 16'h2222;
    PFUMX i23567 (.BLUT(n31670), .ALUT(n31669), .C0(\register_addr[1] ), 
          .Z(n31671));
    PFUMX i23564 (.BLUT(n31667), .ALUT(n31666), .C0(\register_addr[1] ), 
          .Z(n31668));
    LUT4 Select_4249_i2_2_lut (.A(read_value[5]), .B(n52), .Z(n2_adj_444)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4249_i2_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_430 (.A(read_value_adj_264[5]), .B(\read_value[5]_adj_233 ), 
         .C(n46), .D(n31944), .Z(n14_adj_447)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_430.init = 16'heca0;
    LUT4 i2_4_lut_adj_431 (.A(\read_value[5]_adj_234 ), .B(read_value_adj_529[5]), 
         .C(n31942), .D(n46_adj_295), .Z(n12_adj_450)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_431.init = 16'heca0;
    LUT4 i15556_1_lut_4_lut (.A(\register_addr[2] ), .B(n32004), .C(\register_addr[0] ), 
         .D(\register_addr[1] ), .Z(n176)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B))) */ ;
    defparam i15556_1_lut_4_lut.init = 16'h1333;
    L6MUX21 i23527 (.D0(n31590), .D1(n31587), .SD(\register_addr[2] ), 
            .Z(n31591));
    LUT4 i9_4_lut_adj_432 (.A(n17_adj_456), .B(n6_adj_457), .C(n16_adj_458), 
         .D(n2_adj_459), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_432.init = 16'hfffe;
    LUT4 i7_4_lut_adj_433 (.A(\read_value[4]_adj_235 ), .B(n14_adj_461), 
         .C(n5_adj_236), .D(n31924), .Z(n17_adj_456)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_433.init = 16'hfefc;
    PFUMX i23525 (.BLUT(n31589), .ALUT(n31588), .C0(\register_addr[1] ), 
          .Z(n31590));
    PFUMX i23307 (.BLUT(n31007), .ALUT(n31006), .C0(\register_addr[1] ), 
          .Z(n31008));
    FD1S3IX read_value__i0 (.D(n31827), .CK(\select[7] ), .CD(n31949), 
            .Q(read_value_adj_529[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=699, LSE_RLINE=711 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 Select_4250_i6_2_lut (.A(databus_out[4]), .B(n33683), .Z(n6_adj_457)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4250_i6_2_lut.init = 16'h2222;
    LUT4 i9_4_lut_adj_434 (.A(n1), .B(n18), .C(n14_adj_463), .D(n5_adj_237), 
         .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_434.init = 16'hfffe;
    LUT4 i8_4_lut (.A(read_value_adj_264[1]), .B(n16_adj_436), .C(n2_adj_440), 
         .D(n46), .Z(n18)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut.init = 16'hfefc;
    LUT4 i6_4_lut_adj_435 (.A(read_value_adj_265[4]), .B(n12_adj_467), .C(n8_adj_238), 
         .D(n47), .Z(n16_adj_458)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_435.init = 16'hfefc;
    LUT4 Select_4250_i2_2_lut (.A(read_value[4]), .B(n52), .Z(n2_adj_459)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4250_i2_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_436 (.A(read_value_adj_264[4]), .B(\read_value[4]_adj_239 ), 
         .C(n46), .D(n31944), .Z(n14_adj_461)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_436.init = 16'heca0;
    PFUMX i23522 (.BLUT(n31586), .ALUT(n31585), .C0(\register_addr[1] ), 
          .Z(n31587));
    LUT4 i15555_4_lut_rep_332 (.A(\register_addr[2] ), .B(n32004), .C(\register_addr[0] ), 
         .D(\register_addr[1] ), .Z(n31949)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i15555_4_lut_rep_332.init = 16'heccc;
    LUT4 i2_4_lut_adj_437 (.A(\read_value[4]_adj_240 ), .B(read_value_adj_529[4]), 
         .C(n31942), .D(n46_adj_295), .Z(n12_adj_467)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_437.init = 16'heca0;
    L6MUX21 i23496 (.D0(n31529), .D1(n31526), .SD(\register_addr[2] ), 
            .Z(n31530));
    LUT4 i9_4_lut_adj_438 (.A(n17_adj_473), .B(n6_adj_474), .C(n16_adj_475), 
         .D(n2_adj_476), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_438.init = 16'hfffe;
    LUT4 i7_4_lut_adj_439 (.A(\read_value[3]_adj_241 ), .B(n14_adj_478), 
         .C(n5_adj_242), .D(n31924), .Z(n17_adj_473)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_439.init = 16'hfefc;
    PFUMX i23491 (.BLUT(n31525), .ALUT(n31524), .C0(\register_addr[1] ), 
          .Z(n31526));
    LUT4 Select_4251_i6_2_lut (.A(databus_out[3]), .B(rw), .Z(n6_adj_474)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4251_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_440 (.A(read_value_adj_265[3]), .B(n12_adj_481), .C(n8_adj_243), 
         .D(n47), .Z(n16_adj_475)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_440.init = 16'hfefc;
    LUT4 Select_4251_i2_2_lut (.A(read_value[3]), .B(n52), .Z(n2_adj_476)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4251_i2_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_441 (.A(read_value_adj_264[3]), .B(\read_value[3]_adj_244 ), 
         .C(n46), .D(n31944), .Z(n14_adj_478)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_441.init = 16'heca0;
    PFUMX i23494 (.BLUT(n31528), .ALUT(n31527), .C0(\register_addr[1] ), 
          .Z(n31529));
    LUT4 i2_4_lut_adj_442 (.A(\read_value[3]_adj_245 ), .B(read_value_adj_529[3]), 
         .C(n31942), .D(n46_adj_295), .Z(n12_adj_481)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_442.init = 16'heca0;
    LUT4 i9_4_lut_adj_443 (.A(n17_adj_487), .B(n6_adj_488), .C(n16_adj_489), 
         .D(n2_adj_490), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_443.init = 16'hfffe;
    LUT4 i7_4_lut_adj_444 (.A(\read_value[2]_adj_246 ), .B(n14_adj_492), 
         .C(n5_adj_247), .D(n31924), .Z(n17_adj_487)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_444.init = 16'hfefc;
    L6MUX21 i23309 (.D0(n31008), .D1(n31005), .SD(\register_addr[2] ), 
            .Z(n31009));
    LUT4 i4_4_lut_adj_445 (.A(read_value_adj_265[1]), .B(\read_value[1]_adj_248 ), 
         .C(n47), .D(n31944), .Z(n14_adj_463)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_445.init = 16'heca0;
    LUT4 Select_4252_i6_2_lut (.A(databus_out[2]), .B(rw), .Z(n6_adj_488)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4252_i6_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_446 (.A(n9_adj_496), .B(n14_adj_497), .C(n3_adj_249), 
         .D(n5_adj_499), .Z(databus[31])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_446.init = 16'hfffe;
    LUT4 i1_4_lut_adj_447 (.A(\read_value[31]_adj_250 ), .B(read_value_adj_265[31]), 
         .C(n31924), .D(n47), .Z(n9_adj_496)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_447.init = 16'heca0;
    LUT4 i6_4_lut_adj_448 (.A(\read_value[31]_adj_251 ), .B(n12_adj_502), 
         .C(n6_adj_252), .D(n31942), .Z(n14_adj_497)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_448.init = 16'hfefc;
    LUT4 i6_4_lut_adj_449 (.A(read_value_adj_265[2]), .B(n12_adj_505), .C(n8_adj_253), 
         .D(n47), .Z(n16_adj_489)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_449.init = 16'hfefc;
    LUT4 Select_4252_i2_2_lut (.A(read_value[2]), .B(n52), .Z(n2_adj_490)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4252_i2_2_lut.init = 16'h8888;
    LUT4 i9_4_lut_adj_450 (.A(n17_adj_508), .B(n6_adj_509), .C(n16_adj_510), 
         .D(n2_adj_511), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_450.init = 16'hfffe;
    LUT4 i4_4_lut_adj_451 (.A(read_value_adj_264[2]), .B(\read_value[2]_adj_254 ), 
         .C(n46), .D(n31944), .Z(n14_adj_492)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_451.init = 16'heca0;
    LUT4 i7_4_lut_adj_452 (.A(\read_value[0]_adj_255 ), .B(n14_adj_284), 
         .C(n5_adj_256), .D(n31924), .Z(n17_adj_508)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_452.init = 16'hfefc;
    LUT4 Select_4177_i5_2_lut (.A(databus_out[31]), .B(rw), .Z(n5_adj_499)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4177_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_453 (.A(read_value[31]), .B(read_value_adj_264[31]), 
         .C(n52), .D(n46), .Z(n12_adj_502)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_453.init = 16'heca0;
    LUT4 i2_4_lut_adj_454 (.A(\read_value[2]_adj_257 ), .B(read_value_adj_529[2]), 
         .C(n31942), .D(n46_adj_295), .Z(n12_adj_505)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_454.init = 16'heca0;
    LUT4 Select_4254_i6_2_lut (.A(databus_out[0]), .B(rw), .Z(n6_adj_509)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4254_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_455 (.A(read_value_adj_265[0]), .B(n12_adj_296), .C(n8_adj_258), 
         .D(n47), .Z(n16_adj_510)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_455.init = 16'hfefc;
    LUT4 Select_4254_i2_2_lut (.A(read_value[0]), .B(n52), .Z(n2_adj_511)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4254_i2_2_lut.init = 16'h8888;
    PFUMX i23305 (.BLUT(n31004), .ALUT(n31003), .C0(\register_addr[1] ), 
          .Z(n31005));
    PWMReceiver recv_ch8 (.n32039(n32039), .n5(n5_adj_259), .n27979(n27979), 
            .GND_net(GND_net), .debug_c_c(debug_c_c), .n33686(n33686), 
            .rc_ch8_c(rc_ch8_c), .n30381(n30381), .n33685(n33685), .\register[6] ({\register[6] }), 
            .n13735(n13735), .n1234(n1234), .n27956(n27956), .n27877(n27877)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(257[14] 261[36])
    PWMReceiver_U1 recv_ch7 (.debug_c_c(debug_c_c), .n33686(n33686), .rc_ch7_c(rc_ch7_c), 
            .GND_net(GND_net), .n5(n5_adj_260), .n32074(n32074), .n28044(n28044), 
            .n27887(n27887), .n1219(n1219), .n27759(n27759), .n33687(n33687), 
            .\register[5] ({\register[5] }), .n14315(n14315), .n30505(n30505), 
            .n33685(n33685)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(252[14] 256[36])
    PWMReceiver_U2 recv_ch4 (.count({Open_9, Open_10, Open_11, Open_12, 
            Open_13, Open_14, Open_15, \count[8] , Open_16, Open_17, 
            Open_18, Open_19, Open_20, Open_21, Open_22, Open_23}), 
            .GND_net(GND_net), .\count[13] (\count[13] ), .n27644(n27644), 
            .debug_c_c(debug_c_c), .n33686(n33686), .rc_ch4_c(rc_ch4_c), 
            .\count[11] (\count[11] ), .n30520(n30520), .\count[9] (\count[9] ), 
            .\count[10] (\count[10] ), .n32025(n32025), .n154(n154), .n33685(n33685), 
            .n1204(n1204), .n27883(n27883), .n29469(n29469), .n33687(n33687), 
            .\register[4] ({\register[4] }), .n30220(n30220)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(247[14] 251[36])
    PWMReceiver_U3 recv_ch3 (.n5(n5_adj_261), .GND_net(GND_net), .n27879(n27879), 
            .n30196(n30196), .n27809(n27809), .\count[8] (\count[8]_adj_262 ), 
            .n30202(n30202), .\count[9] (\count[9]_adj_263 ), .\count[6] (\count[6] ), 
            .\count[7] (\count[7] ), .n32062(n32062), .\count[5] (\count[5] ), 
            .n27853(n27853), .n32064(n32064), .n27983(n27983), .debug_c_c(debug_c_c), 
            .n33686(n33686), .rc_ch3_c(rc_ch3_c), .n32080(n32080), .n1189(n1189), 
            .n27758(n27758), .n29341(n29341), .n33687(n33687), .\register[3] ({\register[3] }), 
            .n14358(n14358), .n30445(n30445), .n33685(n33685)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(242[14] 246[36])
    PWMReceiver_U4 recv_ch2 (.n1168(n1168), .n1180(n1180), .n31964(n31964), 
            .GND_net(GND_net), .n30426(n30426), .debug_c_c(debug_c_c), 
            .n31906(n31906), .n33687(n33687), .\register[2] ({\register[2] }), 
            .n14369(n14369), .n1174(n1174), .n27757(n27757), .n33685(n33685), 
            .n33686(n33686), .rc_ch2_c(rc_ch2_c), .n29866(n29866)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(237[14] 241[36])
    PWMReceiver_U5 recv_ch1 (.GND_net(GND_net), .n1153(n1153), .debug_c_c(debug_c_c), 
            .n33686(n33686), .n1165(n1165), .n31948(n31948), .n30378(n30378), 
            .\register[1] ({\register[1] }), .n14374(n14374), .n33685(n33685), 
            .rc_ch1_c(rc_ch1_c), .n1159(n1159), .n27960(n27960), .n29869(n29869)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(232[17] 236[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (n32039, n5, n27979, GND_net, debug_c_c, n33686, 
            rc_ch8_c, n30381, n33685, \register[6] , n13735, n1234, 
            n27956, n27877) /* synthesis syn_module_defined=1 */ ;
    output n32039;
    output n5;
    output n27979;
    input GND_net;
    input debug_c_c;
    input n33686;
    input rc_ch8_c;
    output n30381;
    input n33685;
    output [7:0]\register[6] ;
    input n13735;
    output n1234;
    input n27956;
    output n27877;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n32036, n29895, n32037, n30194, n30242, n13527, n31961, 
        n32009, n31993, n32038, n111, n4, n4_adj_165, n29936, 
        n26762;
    wire [15:0]n116;
    
    wire n26763, n1240, n1228, n32058, n32019, n29839, n27703, 
        n31929, n31992, n31963, n27041;
    wire [7:0]n1132;
    
    wire n27040, n29935, n27039, n27038, n54, n29952, n10, n29655, 
        n16775, n26, n30228, n30206;
    wire [7:0]n43;
    
    wire n29896, n26769, n26768, n30159, n26767, n26766, n29627, 
        n26765, n26764;
    
    LUT4 i1_2_lut_rep_419 (.A(count[6]), .B(count[7]), .Z(n32036)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_419.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n29895)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_420 (.A(count[11]), .B(count[10]), .Z(n32037)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_420.init = 16'heeee;
    LUT4 i22786_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[12]), 
         .D(count[13]), .Z(n30194)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22786_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_344_4_lut (.A(count[11]), .B(count[10]), .C(n30242), 
         .D(n13527), .Z(n31961)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_344_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_392_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n32009)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_392_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_376_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n13527), 
         .D(count[9]), .Z(n31993)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_376_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_421 (.A(count[2]), .B(count[1]), .Z(n32038)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_421.init = 16'h8888;
    LUT4 i105_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[3]), .Z(n111)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i105_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_314 (.A(count[2]), .B(count[1]), .C(count[0]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_314.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_315 (.A(count[2]), .B(count[1]), .C(count[4]), 
         .Z(n4_adj_165)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_315.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_422 (.A(count[15]), .B(count[14]), .Z(n32039)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_422.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n27979), 
         .Z(n29936)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n13527)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_1778_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26762), 
          .COUT(n26763), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_3.INIT0 = 16'hd222;
    defparam add_1778_3.INIT1 = 16'hd222;
    defparam add_1778_3.INJECT1_0 = "NO";
    defparam add_1778_3.INJECT1_1 = "NO";
    CCU2D add_1778_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29936), .B1(n1240), .C1(count[0]), .D1(n1228), .COUT(n26762), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_1.INIT0 = 16'hF000;
    defparam add_1778_1.INIT1 = 16'ha565;
    defparam add_1778_1.INJECT1_0 = "NO";
    defparam add_1778_1.INJECT1_1 = "NO";
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n33686), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1240));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1240), .SP(n33686), .CK(debug_c_c), .Q(n1228));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_441 (.A(count[4]), .B(count[5]), .Z(n32058)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_441.init = 16'h8888;
    LUT4 i1_2_lut_rep_402_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n32019)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_402_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_4_lut (.A(n32038), .B(n32036), .C(n32019), .D(count[0]), 
         .Z(n29839)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_312_3_lut_4_lut (.A(n13527), .B(n32009), .C(n27703), 
         .D(count[8]), .Z(n31929)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_312_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_346_4_lut (.A(n13527), .B(n32009), .C(n31992), .D(count[8]), 
         .Z(n31963)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i2_3_lut_rep_346_4_lut.init = 16'hfeff;
    CCU2D sub_79_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27041), 
          .S0(n1132[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_9.INIT1 = 16'h0000;
    defparam sub_79_add_2_9.INJECT1_0 = "NO";
    defparam sub_79_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27040), 
          .COUT(n27041), .S0(n1132[5]), .S1(n1132[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_79_add_2_7.INJECT1_0 = "NO";
    defparam sub_79_add_2_7.INJECT1_1 = "NO";
    LUT4 i23042_3_lut_3_lut_4_lut (.A(n32039), .B(n27979), .C(n31929), 
         .D(n31961), .Z(n29935)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i23042_3_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D sub_79_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27039), 
          .COUT(n27040), .S0(n1132[3]), .S1(n1132[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_79_add_2_5.INJECT1_0 = "NO";
    defparam sub_79_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27038), 
          .COUT(n27039), .S0(n1132[1]), .S1(n1132[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_79_add_2_3.INJECT1_0 = "NO";
    defparam sub_79_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27038), 
          .S1(n1132[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_1.INIT0 = 16'hF000;
    defparam sub_79_add_2_1.INIT1 = 16'h5555;
    defparam sub_79_add_2_1.INJECT1_0 = "NO";
    defparam sub_79_add_2_1.INJECT1_1 = "NO";
    LUT4 i3_3_lut_rep_375_4_lut (.A(count[3]), .B(n32058), .C(n32036), 
         .D(n32038), .Z(n31992)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_3_lut_rep_375_4_lut.init = 16'h8000;
    LUT4 i23069_4_lut (.A(n54), .B(n29952), .C(n31963), .D(n10), .Z(n30381)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23069_4_lut.init = 16'h3323;
    LUT4 i3_4_lut (.A(n32039), .B(n29655), .C(n30242), .D(n33685), .Z(n16775)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i6_4_lut (.A(n26), .B(n30194), .C(n1228), .D(n1240), .Z(n29655)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i6_4_lut.init = 16'h0020;
    LUT4 i1_4_lut (.A(n29895), .B(n31993), .C(n32019), .D(n4), .Z(n26)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut.init = 16'heccc;
    LUT4 i22834_3_lut (.A(count[9]), .B(count[8]), .C(n30228), .Z(n30242)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i22834_3_lut.init = 16'ha8a8;
    LUT4 i22820_4_lut (.A(n30206), .B(count[7]), .C(n32058), .D(count[6]), 
         .Z(n30228)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;
    defparam i22820_4_lut.init = 16'hffec;
    LUT4 i22798_4_lut (.A(count[3]), .B(count[1]), .C(count[2]), .D(count[0]), 
         .Z(n30206)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22798_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n32036), .B(count[5]), .C(count[3]), .D(n4_adj_165), 
         .Z(n27703)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_2_lut (.A(n1240), .B(n1228), .Z(n29952)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i5_2_lut (.A(n1228), .B(n1240), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_316 (.A(count[13]), .B(count[12]), .C(n29896), .D(n32009), 
         .Z(n27979)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_316.init = 16'h8880;
    CCU2D add_1778_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26769), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_17.INIT0 = 16'hd222;
    defparam add_1778_17.INIT1 = 16'h0000;
    defparam add_1778_17.INJECT1_0 = "NO";
    defparam add_1778_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_317 (.A(count[4]), .B(n29895), .C(n111), .D(count[5]), 
         .Z(n29896)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_317.init = 16'hccc8;
    CCU2D add_1778_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26768), 
          .COUT(n26769), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_15.INIT0 = 16'hd222;
    defparam add_1778_15.INIT1 = 16'hd222;
    defparam add_1778_15.INJECT1_0 = "NO";
    defparam add_1778_15.INJECT1_1 = "NO";
    LUT4 i21_2_lut_4_lut (.A(n13527), .B(n30242), .C(n32037), .D(n26), 
         .Z(n54)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i21_2_lut_4_lut.init = 16'h0100;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31993), .C(n29839), 
         .D(n27703), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(160[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22751_3_lut_4_lut (.A(count[8]), .B(n31993), .C(n27703), .D(n29839), 
         .Z(n30159)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(160[28:39])
    defparam i22751_3_lut_4_lut.init = 16'hfeee;
    CCU2D add_1778_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26767), 
          .COUT(n26768), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_13.INIT0 = 16'hd222;
    defparam add_1778_13.INIT1 = 16'hd222;
    defparam add_1778_13.INJECT1_0 = "NO";
    defparam add_1778_13.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13735), .PD(n16775), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1778_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26766), 
          .COUT(n26767), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_11.INIT0 = 16'hd222;
    defparam add_1778_11.INIT1 = 16'hd222;
    defparam add_1778_11.INJECT1_0 = "NO";
    defparam add_1778_11.INJECT1_1 = "NO";
    LUT4 i15390_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15390_2_lut_4_lut.init = 16'h0400;
    LUT4 i15389_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15389_2_lut_4_lut.init = 16'h0400;
    LUT4 i15388_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15388_2_lut_4_lut.init = 16'h0400;
    LUT4 i15387_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15387_2_lut_4_lut.init = 16'h0400;
    LUT4 i15386_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15386_2_lut_4_lut.init = 16'h0400;
    LUT4 i15385_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15385_2_lut_4_lut.init = 16'h0400;
    LUT4 i15384_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15384_2_lut_4_lut.init = 16'h0400;
    LUT4 i15134_2_lut_4_lut (.A(n31993), .B(count[8]), .C(n31992), .D(n1132[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15134_2_lut_4_lut.init = 16'h0400;
    FD1P3AX valid_48 (.D(n29935), .SP(n27956), .CK(debug_c_c), .Q(n1234));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_318 (.A(n30159), .B(n29952), .C(n30242), .D(n29627), 
         .Z(n27877)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_318.init = 16'hcecc;
    LUT4 i3_4_lut_adj_319 (.A(n54), .B(n32037), .C(n31963), .D(n13527), 
         .Z(n29627)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_319.init = 16'h0010;
    CCU2D add_1778_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26765), 
          .COUT(n26766), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_9.INIT0 = 16'hd222;
    defparam add_1778_9.INIT1 = 16'hd222;
    defparam add_1778_9.INJECT1_0 = "NO";
    defparam add_1778_9.INJECT1_1 = "NO";
    CCU2D add_1778_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26764), 
          .COUT(n26765), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_7.INIT0 = 16'hd222;
    defparam add_1778_7.INIT1 = 16'hd222;
    defparam add_1778_7.INJECT1_0 = "NO";
    defparam add_1778_7.INJECT1_1 = "NO";
    CCU2D add_1778_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26763), 
          .COUT(n26764), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1778_5.INIT0 = 16'hd222;
    defparam add_1778_5.INIT1 = 16'hd222;
    defparam add_1778_5.INJECT1_0 = "NO";
    defparam add_1778_5.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (debug_c_c, n33686, rc_ch7_c, GND_net, n5, n32074, 
            n28044, n27887, n1219, n27759, n33687, \register[5] , 
            n14315, n30505, n33685) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n33686;
    input rc_ch7_c;
    input GND_net;
    output n5;
    output n32074;
    output n28044;
    output n27887;
    output n1219;
    input n27759;
    input n33687;
    output [7:0]\register[5] ;
    input n14315;
    output n30505;
    input n33685;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27634, n31974, n33678, n31939, n29986, n27767, n13424;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n10, n31973;
    wire [7:0]n1123;
    
    wire n29602;
    wire [7:0]n43;
    
    wire n1213, n1225, n31997, n32069, n29429, n32070, n32023, 
        n32071, n32022, n4, n27045, n27044, n26777;
    wire [15:0]n116;
    
    wire n26776, n27043, n4_adj_161, n27042, n32073, n30198, n29987, 
        n5_adj_162, n30120, n30147, n26775, n27923, n6, n29751, 
        n4_adj_163, n26774, n26773, n26772, n16596, n26771, n26770, 
        n10_adj_164, n11;
    
    LUT4 i23180_3_lut_3_lut_4_lut (.A(n27634), .B(n31974), .C(n33678), 
         .D(n31939), .Z(n29986)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23180_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i15665_3_lut_rep_474 (.A(n27767), .B(n13424), .C(count[9]), .Z(n33678)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15665_3_lut_rep_474.init = 16'hecec;
    LUT4 i21_3_lut_rep_356_4_lut_4_lut (.A(n27767), .B(n13424), .C(count[9]), 
         .D(n10), .Z(n31973)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i21_3_lut_rep_356_4_lut_4_lut.init = 16'h1310;
    LUT4 i15375_2_lut (.A(n1123[1]), .B(n29602), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15375_2_lut.init = 16'h2222;
    FD1P3AX prev_in_46 (.D(n1225), .SP(n33686), .CK(debug_c_c), .Q(n1213));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n33686), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1225));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_380 (.A(count[9]), .B(n13424), .Z(n31997)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_380.init = 16'heeee;
    LUT4 i1_2_lut_rep_357_3_lut (.A(count[9]), .B(n13424), .C(count[8]), 
         .Z(n31974)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_357_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_452 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n32069)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_452.init = 16'h8080;
    LUT4 i1_2_lut_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), .D(count[0]), 
         .Z(n29429)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i14917_2_lut_rep_453 (.A(count[5]), .B(count[4]), .Z(n32070)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14917_2_lut_rep_453.init = 16'h8888;
    LUT4 i2_3_lut_rep_406_4_lut (.A(count[5]), .B(count[4]), .C(count[6]), 
         .D(count[7]), .Z(n32023)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_406_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_454 (.A(count[6]), .B(count[7]), .Z(n32071)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_454.init = 16'h8888;
    LUT4 i1_2_lut_rep_405_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n32022)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_405_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    CCU2D sub_78_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27045), 
          .S0(n1123[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_9.INIT1 = 16'h0000;
    defparam sub_78_add_2_9.INJECT1_0 = "NO";
    defparam sub_78_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27044), 
          .COUT(n27045), .S0(n1123[5]), .S1(n1123[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_7.INJECT1_0 = "NO";
    defparam sub_78_add_2_7.INJECT1_1 = "NO";
    CCU2D add_1774_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26777), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_17.INIT0 = 16'hd222;
    defparam add_1774_17.INIT1 = 16'h0000;
    defparam add_1774_17.INJECT1_0 = "NO";
    defparam add_1774_17.INJECT1_1 = "NO";
    CCU2D add_1774_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26776), 
          .COUT(n26777), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_15.INIT0 = 16'hd222;
    defparam add_1774_15.INIT1 = 16'hd222;
    defparam add_1774_15.INJECT1_0 = "NO";
    defparam add_1774_15.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27043), 
          .COUT(n27044), .S0(n1123[3]), .S1(n1123[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_5.INJECT1_0 = "NO";
    defparam sub_78_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_161)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    CCU2D sub_78_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27042), 
          .COUT(n27043), .S0(n1123[1]), .S1(n1123[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_3.INJECT1_0 = "NO";
    defparam sub_78_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_456 (.A(count[11]), .B(count[10]), .Z(n32073)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_456.init = 16'heeee;
    LUT4 i22790_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n30198)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22790_3_lut_4_lut.init = 16'hfffe;
    CCU2D sub_78_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27042), 
          .S1(n1123[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_1.INIT0 = 16'hF000;
    defparam sub_78_add_2_1.INIT1 = 16'h5555;
    defparam sub_78_add_2_1.INJECT1_0 = "NO";
    defparam sub_78_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_457 (.A(count[15]), .B(count[14]), .Z(n32074)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_457.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n28044), 
         .Z(n29987)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_322_3_lut (.A(count[15]), .B(count[14]), .C(n28044), 
         .Z(n31939)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_322_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut (.A(n5_adj_162), .B(n30120), .C(n30147), .D(n33678), 
         .Z(n27887)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    CCU2D add_1774_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26775), 
          .COUT(n26776), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_13.INIT0 = 16'hd222;
    defparam add_1774_13.INIT1 = 16'hd222;
    defparam add_1774_13.INJECT1_0 = "NO";
    defparam add_1774_13.INJECT1_1 = "NO";
    LUT4 i3_4_lut (.A(n27923), .B(n6), .C(count[8]), .D(n32070), .Z(n27767)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut.init = 16'hfefc;
    LUT4 i3_4_lut_adj_306 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27923)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_306.init = 16'hfffe;
    LUT4 i5_2_lut (.A(n1213), .B(n1225), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_307 (.A(count[12]), .B(count[13]), .C(n32074), .D(n32073), 
         .Z(n13424)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_307.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n32071), .B(count[4]), .C(count[5]), .D(n4), .Z(n27634)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i3_3_lut_4_lut (.A(count[8]), .B(n32071), .C(n29429), .D(n32070), 
         .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_308 (.A(count[7]), .B(count[6]), .C(n32070), 
         .D(n29429), .Z(n29751)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_308.init = 16'h8000;
    FD1P3AX valid_48 (.D(n29986), .SP(n27759), .CK(debug_c_c), .Q(n1219));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_309 (.A(n31997), .B(count[8]), .C(n32023), .D(n32069), 
         .Z(n29602)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_309.init = 16'hfbbb;
    LUT4 i22716_2_lut (.A(n1213), .B(n1225), .Z(n30120)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22716_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_adj_310 (.A(count[13]), .B(count[12]), .C(n32073), .D(n4_adj_163), 
         .Z(n28044)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_310.init = 16'h8880;
    LUT4 i1_4_lut_adj_311 (.A(count[5]), .B(count[9]), .C(n32022), .D(n4_adj_161), 
         .Z(n4_adj_163)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_311.init = 16'hfcec;
    CCU2D add_1774_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26774), 
          .COUT(n26775), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_11.INIT0 = 16'hd222;
    defparam add_1774_11.INIT1 = 16'hd222;
    defparam add_1774_11.INJECT1_0 = "NO";
    defparam add_1774_11.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    CCU2D add_1774_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26773), 
          .COUT(n26774), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_9.INIT0 = 16'hd222;
    defparam add_1774_9.INIT1 = 16'hd222;
    defparam add_1774_9.INJECT1_0 = "NO";
    defparam add_1774_9.INJECT1_1 = "NO";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    CCU2D add_1774_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26772), 
          .COUT(n26773), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_7.INIT0 = 16'hd222;
    defparam add_1774_7.INIT1 = 16'hd222;
    defparam add_1774_7.INJECT1_0 = "NO";
    defparam add_1774_7.INJECT1_1 = "NO";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    CCU2D add_1774_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26771), 
          .COUT(n26772), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_5.INIT0 = 16'hd222;
    defparam add_1774_5.INIT1 = 16'hd222;
    defparam add_1774_5.INJECT1_0 = "NO";
    defparam add_1774_5.INJECT1_1 = "NO";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1774_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26770), 
          .COUT(n26771), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_3.INIT0 = 16'hd222;
    defparam add_1774_3.INIT1 = 16'hd222;
    defparam add_1774_3.INJECT1_0 = "NO";
    defparam add_1774_3.INJECT1_1 = "NO";
    CCU2D add_1774_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29987), .B1(n1225), .C1(count[0]), .D1(n1213), .COUT(n26770), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1774_1.INIT0 = 16'hF000;
    defparam add_1774_1.INIT1 = 16'ha565;
    defparam add_1774_1.INJECT1_0 = "NO";
    defparam add_1774_1.INJECT1_1 = "NO";
    LUT4 i15378_2_lut (.A(n1123[4]), .B(n29602), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15378_2_lut.init = 16'h2222;
    LUT4 i15377_2_lut (.A(n1123[3]), .B(n29602), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15377_2_lut.init = 16'h2222;
    LUT4 i15379_2_lut (.A(n1123[5]), .B(n29602), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15379_2_lut.init = 16'h2222;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14315), .PD(n16596), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i15129_2_lut (.A(n1123[0]), .B(n29602), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15129_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_4_lut_adj_312 (.A(n10), .B(n33678), .C(n31997), .D(n29602), 
         .Z(n5_adj_162)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut_adj_312.init = 16'hcd00;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31997), .C(n29751), 
         .D(n27634), .Z(n10_adj_164)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(160[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22742_3_lut_4_lut (.A(count[8]), .B(n31997), .C(n27634), .D(n29751), 
         .Z(n30147)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(160[28:39])
    defparam i22742_3_lut_4_lut.init = 16'hfeee;
    LUT4 i23193_4_lut (.A(n31973), .B(n30120), .C(n29602), .D(n10_adj_164), 
         .Z(n30505)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23193_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_313 (.A(n33685), .B(n32074), .C(n11), .D(n30198), 
         .Z(n16596)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_313.init = 16'h0020;
    LUT4 i4_4_lut (.A(n10), .B(n30120), .C(n27767), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i15381_2_lut (.A(n1123[7]), .B(n29602), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15381_2_lut.init = 16'h2222;
    LUT4 i15376_2_lut (.A(n1123[2]), .B(n29602), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15376_2_lut.init = 16'h2222;
    LUT4 i15380_2_lut (.A(n1123[6]), .B(n29602), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15380_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (count, GND_net, \count[13] , n27644, debug_c_c, 
            n33686, rc_ch4_c, \count[11] , n30520, \count[9] , \count[10] , 
            n32025, n154, n33685, n1204, n27883, n29469, n33687, 
            \register[4] , n30220) /* synthesis syn_module_defined=1 */ ;
    output [15:0]count;
    input GND_net;
    output \count[13] ;
    output n27644;
    input debug_c_c;
    input n33686;
    input rc_ch4_c;
    output \count[11] ;
    output n30520;
    output \count[9] ;
    output \count[10] ;
    output n32025;
    output n154;
    input n33685;
    output n1204;
    input n27883;
    input n29469;
    input n33687;
    output [7:0]\register[4] ;
    input n30220;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n31976, n31999, n54, n5;
    wire [7:0]n1114;
    wire [7:0]n43;
    
    wire n1198, n1210, n32040, n28045, n32085, n28074, n26785;
    wire [15:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    wire [15:0]n116;
    
    wire n26784, n29756, n30149, n26783, n27882, n32076, n30046, 
        n26782, n32083, n4, n26781, n32091, n32092, n32093, n31998, 
        n5_adj_157, n6, n29973, n32084, n32024, n26780, n26779, 
        n27049, n27048, n26778, n27047, n27046, n4_adj_158, n32072, 
        n32077, n103, n32031, n4_adj_159, n14349, n6_adj_160, n152, 
        n16629, n26;
    
    LUT4 i1_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n54), 
         .Z(n5)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h00fb;
    LUT4 i15374_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15374_2_lut_4_lut.init = 16'h0400;
    LUT4 i5_2_lut_rep_423 (.A(n1198), .B(n1210), .Z(n32040)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_423.init = 16'h4444;
    LUT4 i15373_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15373_2_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_4_lut (.A(n1198), .B(n1210), .C(n28045), .D(n32085), 
         .Z(n28074)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i2_3_lut_4_lut.init = 16'hfff4;
    LUT4 i15372_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15372_2_lut_4_lut.init = 16'h0400;
    LUT4 i15371_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15371_2_lut_4_lut.init = 16'h0400;
    LUT4 i15370_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15370_2_lut_4_lut.init = 16'h0400;
    CCU2D add_1770_17 (.A0(count_c[15]), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26785), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_17.INIT0 = 16'hd222;
    defparam add_1770_17.INIT1 = 16'h0000;
    defparam add_1770_17.INJECT1_0 = "NO";
    defparam add_1770_17.INJECT1_1 = "NO";
    LUT4 i15369_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15369_2_lut_4_lut.init = 16'h0400;
    CCU2D add_1770_15 (.A0(\count[13] ), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[14]), .B1(n32040), .C1(GND_net), .D1(GND_net), 
          .CIN(n26784), .COUT(n26785), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_15.INIT0 = 16'hd222;
    defparam add_1770_15.INIT1 = 16'hd222;
    defparam add_1770_15.INJECT1_0 = "NO";
    defparam add_1770_15.INJECT1_1 = "NO";
    LUT4 i15368_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15368_2_lut_4_lut.init = 16'h0400;
    LUT4 i15124_2_lut_4_lut (.A(n31976), .B(count[8]), .C(n31999), .D(n1114[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15124_2_lut_4_lut.init = 16'h0400;
    LUT4 i22743_3_lut_4_lut (.A(count[8]), .B(n31976), .C(n27644), .D(n29756), 
         .Z(n30149)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22743_3_lut_4_lut.init = 16'hfeee;
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n33686), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1210));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1210), .SP(n33686), .CK(debug_c_c), .Q(n1198));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D add_1770_13 (.A0(\count[11] ), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[12]), .B1(n32040), .C1(GND_net), .D1(GND_net), 
          .CIN(n26783), .COUT(n26784), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_13.INIT0 = 16'hd222;
    defparam add_1770_13.INIT1 = 16'hd222;
    defparam add_1770_13.INJECT1_0 = "NO";
    defparam add_1770_13.INJECT1_1 = "NO";
    LUT4 i23208_4_lut (.A(n32085), .B(n32040), .C(n28045), .D(n27882), 
         .Z(n30520)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23208_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5), .B(n32076), .C(n30149), .D(n30046), .Z(n27882)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    CCU2D add_1770_11 (.A0(\count[9] ), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(\count[10] ), .B1(n32040), .C1(GND_net), .D1(GND_net), 
          .CIN(n26782), .COUT(n26783), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_11.INIT0 = 16'hd222;
    defparam add_1770_11.INIT1 = 16'hd222;
    defparam add_1770_11.INJECT1_0 = "NO";
    defparam add_1770_11.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n32083), .B(count_c[5]), .C(count_c[3]), .D(n4), 
         .Z(n27644)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut.init = 16'h8880;
    CCU2D add_1770_9 (.A0(count_c[7]), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32040), .C1(GND_net), .D1(GND_net), .CIN(n26781), 
          .COUT(n26782), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_9.INIT0 = 16'hd222;
    defparam add_1770_9.INIT1 = 16'hd222;
    defparam add_1770_9.INJECT1_0 = "NO";
    defparam add_1770_9.INJECT1_1 = "NO";
    PFUMX i23662 (.BLUT(n32091), .ALUT(n32092), .C0(count[8]), .Z(n32093));
    LUT4 i1_4_lut_then_3_lut (.A(\count[9] ), .B(n31998), .C(n31999), 
         .Z(n32092)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i1_4_lut_then_3_lut.init = 16'h0101;
    LUT4 i21_4_lut (.A(n5_adj_157), .B(n30046), .C(n31976), .D(n6), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_2_lut_rep_359_4_lut (.A(n32025), .B(\count[13] ), .C(n29973), 
         .D(\count[9] ), .Z(n31976)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_359_4_lut.init = 16'hfffe;
    LUT4 i22644_3_lut (.A(n31998), .B(\count[9] ), .C(n154), .Z(n30046)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i22644_3_lut.init = 16'heaea;
    LUT4 i1_2_lut_4_lut_adj_301 (.A(n32084), .B(n32083), .C(n32024), .D(count_c[0]), 
         .Z(n29756)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_301.init = 16'h8000;
    CCU2D add_1770_7 (.A0(count_c[5]), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[6]), .B1(n32040), .C1(GND_net), .D1(GND_net), 
          .CIN(n26780), .COUT(n26781), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_7.INIT0 = 16'hd222;
    defparam add_1770_7.INIT1 = 16'hd222;
    defparam add_1770_7.INJECT1_0 = "NO";
    defparam add_1770_7.INJECT1_1 = "NO";
    CCU2D add_1770_5 (.A0(count_c[3]), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[4]), .B1(n32040), .C1(GND_net), .D1(GND_net), 
          .CIN(n26779), .COUT(n26780), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_5.INIT0 = 16'hd222;
    defparam add_1770_5.INIT1 = 16'hd222;
    defparam add_1770_5.INJECT1_0 = "NO";
    defparam add_1770_5.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_9 (.A0(count_c[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27049), .S0(n1114[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_9.INIT1 = 16'h0000;
    defparam sub_77_add_2_9.INJECT1_0 = "NO";
    defparam sub_77_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_7 (.A0(count_c[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27048), .COUT(n27049), .S0(n1114[5]), 
          .S1(n1114[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_7.INJECT1_0 = "NO";
    defparam sub_77_add_2_7.INJECT1_1 = "NO";
    CCU2D add_1770_3 (.A0(count_c[1]), .B0(n32040), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[2]), .B1(n32040), .C1(GND_net), .D1(GND_net), 
          .CIN(n26778), .COUT(n26779), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_3.INIT0 = 16'hd222;
    defparam add_1770_3.INIT1 = 16'hd222;
    defparam add_1770_3.INJECT1_0 = "NO";
    defparam add_1770_3.INJECT1_1 = "NO";
    CCU2D add_1770_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28074), .B1(n1210), .C1(count_c[0]), .D1(n1198), .COUT(n26778), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1770_1.INIT0 = 16'hF000;
    defparam add_1770_1.INIT1 = 16'ha565;
    defparam add_1770_1.INJECT1_0 = "NO";
    defparam add_1770_1.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_5 (.A0(count_c[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27047), .COUT(n27048), .S0(n1114[3]), 
          .S1(n1114[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_5.INJECT1_0 = "NO";
    defparam sub_77_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_3 (.A0(count_c[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27046), .COUT(n27047), .S0(n1114[1]), 
          .S1(n1114[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_3.INJECT1_0 = "NO";
    defparam sub_77_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27046), .S1(n1114[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_1.INIT0 = 16'hF000;
    defparam sub_77_add_2_1.INIT1 = 16'h5555;
    defparam sub_77_add_2_1.INJECT1_0 = "NO";
    defparam sub_77_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_302 (.A(\count[13] ), .B(count_c[12]), .C(n29973), 
         .D(n4_adj_158), .Z(n28045)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_302.init = 16'h8880;
    LUT4 i2_3_lut_rep_455 (.A(count_c[7]), .B(count_c[6]), .C(count[8]), 
         .Z(n32072)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_455.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_303 (.A(count_c[7]), .B(count_c[6]), .C(count[8]), 
         .D(n32077), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_303.init = 16'hfffe;
    LUT4 i1_4_lut_adj_304 (.A(\count[9] ), .B(count_c[4]), .C(n32031), 
         .D(n4_adj_159), .Z(n4_adj_158)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_304.init = 16'hfaea;
    LUT4 i1_2_lut (.A(\count[10] ), .B(\count[11] ), .Z(n29973)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i22740_2_lut_rep_459 (.A(n1198), .B(n1210), .Z(n32076)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22740_2_lut_rep_459.init = 16'hdddd;
    LUT4 i1_2_lut_rep_460 (.A(count_c[4]), .B(count_c[5]), .Z(n32077)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_460.init = 16'h8888;
    LUT4 i1_2_lut_rep_407_3_lut (.A(count_c[4]), .B(count_c[5]), .C(count_c[3]), 
         .Z(n32024)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_407_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count_c[4]), .B(count_c[5]), .C(count_c[0]), 
         .D(count_c[3]), .Z(n5_adj_157)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_else_3_lut (.A(\count[9] ), .B(n27644), .C(n29756), 
         .D(n31998), .Z(n32091)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_else_3_lut.init = 16'h0004;
    LUT4 i23192_4_lut_4_lut (.A(n32076), .B(n32093), .C(n33685), .D(n54), 
         .Z(n14349)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23192_4_lut_4_lut.init = 16'h5040;
    LUT4 i23_4_lut (.A(n32072), .B(count_c[2]), .C(n32077), .D(n6_adj_160), 
         .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count_c[1]), .B(count_c[0]), .Z(n6_adj_160)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_466 (.A(count_c[7]), .B(count_c[6]), .Z(n32083)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_466.init = 16'h8888;
    LUT4 i3_3_lut_rep_382_4_lut (.A(count_c[3]), .B(n32077), .C(n32083), 
         .D(n32084), .Z(n31999)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_3_lut_rep_382_4_lut.init = 16'h8000;
    FD1P3AX valid_48 (.D(n29469), .SP(n27883), .CK(debug_c_c), .Q(n1204));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_414_3_lut (.A(count_c[7]), .B(count_c[6]), .C(count[8]), 
         .Z(n32031)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_414_3_lut.init = 16'h8080;
    LUT4 i3_3_lut_rep_381_4_lut (.A(count_c[12]), .B(n32085), .C(n29973), 
         .D(\count[13] ), .Z(n31998)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_381_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count_c[7]), .B(count_c[6]), .C(n32084), 
         .D(count[8]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_467 (.A(count_c[2]), .B(count_c[1]), .Z(n32084)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_467.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(count_c[2]), .B(count_c[1]), .C(count_c[5]), 
         .D(count_c[3]), .Z(n4_adj_159)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_3_lut (.A(count_c[2]), .B(count_c[1]), .C(count_c[4]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_468 (.A(count_c[15]), .B(count_c[14]), .Z(n32085)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_468.init = 16'heeee;
    LUT4 i1_2_lut_rep_408_3_lut (.A(count_c[15]), .B(count_c[14]), .C(count_c[12]), 
         .Z(n32025)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_408_3_lut.init = 16'hfefe;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count_c[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count_c[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[13] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count_c[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[11] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[10] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count_c[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count_c[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count_c[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count_c[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count_c[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count_c[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count_c[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    PFUMX i14223 (.BLUT(n152), .ALUT(n103), .C0(count_c[3]), .Z(n154));
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count_c[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14349), .PD(n16629), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_305 (.A(n33685), .B(n30220), .C(n26), .D(n32076), 
         .Z(n16629)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_305.init = 16'h0020;
    LUT4 i33_4_lut (.A(count[8]), .B(n154), .C(\count[9] ), .D(n29756), 
         .Z(n26)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_4_lut.init = 16'h3a30;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (n5, GND_net, n27879, n30196, n27809, \count[8] , 
            n30202, \count[9] , \count[6] , \count[7] , n32062, \count[5] , 
            n27853, n32064, n27983, debug_c_c, n33686, rc_ch3_c, 
            n32080, n1189, n27758, n29341, n33687, \register[3] , 
            n14358, n30445, n33685) /* synthesis syn_module_defined=1 */ ;
    output n5;
    input GND_net;
    output n27879;
    output n30196;
    output n27809;
    output \count[8] ;
    input n30202;
    output \count[9] ;
    output \count[6] ;
    output \count[7] ;
    output n32062;
    output \count[5] ;
    output n27853;
    output n32064;
    output n27983;
    input debug_c_c;
    input n33686;
    input rc_ch3_c;
    output n32080;
    output n1189;
    input n27758;
    input n29341;
    input n33687;
    output [7:0]\register[3] ;
    input n14358;
    output n30445;
    input n33685;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26787;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    wire [15:0]n116;
    
    wire n26788, n26786, n28072, n1195, n1183, n5_adj_154, n30150, 
        n30153, n33679, n32029, n31978, n32079, n32028, n4, n32027, 
        n32026, n10, n32000, n29746, n29902, n10_adj_155, n31945, 
        n32063, n27053;
    wire [7:0]n1105;
    
    wire n27052, n27051, n27050, n29937, n16639;
    wire [7:0]n43;
    
    wire n4_adj_156, n27895, n26, n26793, n26792, n26791, n26790, 
        n26789;
    
    CCU2D add_1766_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26787), 
          .COUT(n26788), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_5.INIT0 = 16'hd222;
    defparam add_1766_5.INIT1 = 16'hd222;
    defparam add_1766_5.INJECT1_0 = "NO";
    defparam add_1766_5.INJECT1_1 = "NO";
    CCU2D add_1766_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26786), 
          .COUT(n26787), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_3.INIT0 = 16'hd222;
    defparam add_1766_3.INIT1 = 16'hd222;
    defparam add_1766_3.INJECT1_0 = "NO";
    defparam add_1766_3.INJECT1_1 = "NO";
    CCU2D add_1766_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28072), .B1(n1195), .C1(count[0]), .D1(n1183), .COUT(n26786), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_1.INIT0 = 16'hF000;
    defparam add_1766_1.INIT1 = 16'ha565;
    defparam add_1766_1.INJECT1_0 = "NO";
    defparam add_1766_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n5_adj_154), .B(n30150), .C(n30153), .D(n33679), 
         .Z(n27879)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i22788_4_lut (.A(count[13]), .B(count[10]), .C(count[11]), .D(n32029), 
         .Z(n30196)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22788_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27809)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n31978), .B(\count[8] ), .C(n32079), .D(n32028), 
         .Z(n4)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i2_4_lut.init = 16'hfbbb;
    LUT4 i3_4_lut_adj_294 (.A(count[4]), .B(n32027), .C(\count[8] ), .D(n32026), 
         .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_294.init = 16'h8000;
    LUT4 i5_2_lut (.A(n1183), .B(n1195), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i22638_3_lut_rep_475 (.A(n30202), .B(n32000), .C(\count[9] ), 
         .Z(n33679)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i22638_3_lut_rep_475.init = 16'hecec;
    LUT4 i22746_3_lut_4_lut (.A(\count[8] ), .B(n31978), .C(n29746), .D(n29902), 
         .Z(n30153)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22746_3_lut_4_lut.init = 16'hfeee;
    LUT4 i10_3_lut_4_lut (.A(\count[8] ), .B(n31978), .C(n29902), .D(n29746), 
         .Z(n10_adj_155)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_4_lut.init = 16'h0100;
    LUT4 i22744_2_lut (.A(n1183), .B(n1195), .Z(n30150)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22744_2_lut.init = 16'hdddd;
    LUT4 i21_3_lut_rep_328_4_lut_4_lut (.A(n30202), .B(n32000), .C(\count[9] ), 
         .D(n10), .Z(n31945)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i21_3_lut_rep_328_4_lut_4_lut.init = 16'h1310;
    LUT4 i1_2_lut_rep_445 (.A(\count[6] ), .B(\count[7] ), .Z(n32062)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_445.init = 16'h8888;
    LUT4 i1_2_lut_rep_409_3_lut (.A(\count[6] ), .B(\count[7] ), .C(\count[5] ), 
         .Z(n32026)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_409_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\count[6] ), .B(\count[7] ), .C(n27853), 
         .D(\count[5] ), .Z(n29746)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i3145_2_lut_rep_446 (.A(count[1]), .B(count[2]), .Z(n32063)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3145_2_lut_rep_446.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n27853)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_447 (.A(count[15]), .B(count[14]), .Z(n32064)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_447.init = 16'heeee;
    LUT4 i1_2_lut_rep_412_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n32029)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_412_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut_adj_295 (.A(count[15]), .B(count[14]), .C(n5), 
         .D(n27983), .Z(n28072)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_295.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(n10), .B(n33679), .C(n31978), .D(n4), .Z(n5_adj_154)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    CCU2D sub_76_add_2_9 (.A0(\count[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27053), .S0(n1105[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_9.INIT1 = 16'h0000;
    defparam sub_76_add_2_9.INJECT1_0 = "NO";
    defparam sub_76_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27052), .COUT(n27053), .S0(n1105[5]), 
          .S1(n1105[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_7.INJECT1_0 = "NO";
    defparam sub_76_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27051), 
          .COUT(n27052), .S0(n1105[3]), .S1(n1105[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_5.INJECT1_0 = "NO";
    defparam sub_76_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27050), 
          .COUT(n27051), .S0(n1105[1]), .S1(n1105[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_3.INJECT1_0 = "NO";
    defparam sub_76_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27050), 
          .S1(n1105[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_1.INIT0 = 16'hF000;
    defparam sub_76_add_2_1.INIT1 = 16'h5555;
    defparam sub_76_add_2_1.INJECT1_0 = "NO";
    defparam sub_76_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_361_4_lut (.A(n32029), .B(count[13]), .C(n29937), 
         .D(\count[9] ), .Z(n31978)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_361_4_lut.init = 16'hfffe;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n33686), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1195));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_462 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n32079)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_462.init = 16'h8080;
    LUT4 i1_2_lut_rep_410_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n32027)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_410_4_lut.init = 16'h8000;
    LUT4 i14873_2_lut_rep_463 (.A(count[4]), .B(\count[5] ), .Z(n32080)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14873_2_lut_rep_463.init = 16'h8888;
    LUT4 i1_2_lut_rep_411_3_lut_4_lut (.A(count[4]), .B(\count[5] ), .C(\count[7] ), 
         .D(\count[6] ), .Z(n32028)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_411_3_lut_4_lut.init = 16'h8000;
    FD1P3AX valid_48 (.D(n29341), .SP(n27758), .CK(debug_c_c), .Q(n1189));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1195), .SP(n33686), .CK(debug_c_c), .Q(n1183));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_296 (.A(n32080), .B(n32062), .C(n32079), 
         .D(count[0]), .Z(n29902)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_296.init = 16'h8000;
    LUT4 i3_3_lut_rep_383_4_lut (.A(count[12]), .B(n32064), .C(n29937), 
         .D(count[13]), .Z(n32000)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_383_4_lut.init = 16'hfffe;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[7] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_297 (.A(count[13]), .B(count[12]), .C(n29937), .D(n4_adj_156), 
         .Z(n27983)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_297.init = 16'h8880;
    LUT4 i1_4_lut_adj_298 (.A(n32062), .B(\count[9] ), .C(n27895), .D(\count[8] ), 
         .Z(n4_adj_156)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_298.init = 16'heccc;
    LUT4 i2_4_lut_adj_299 (.A(\count[5] ), .B(count[4]), .C(n32063), .D(count[3]), 
         .Z(n27895)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_299.init = 16'hfeee;
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n29937)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i23133_4_lut (.A(n31945), .B(n30150), .C(n4), .D(n10_adj_155), 
         .Z(n30445)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23133_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_300 (.A(n33685), .B(n30196), .C(n26), .D(n30150), 
         .Z(n16639)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_300.init = 16'h0020;
    LUT4 i33_3_lut (.A(n10), .B(n30202), .C(\count[9] ), .Z(n26)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_3_lut.init = 16'h3a3a;
    LUT4 i15363_2_lut (.A(n1105[7]), .B(n4), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15363_2_lut.init = 16'h2222;
    LUT4 i15362_2_lut (.A(n1105[6]), .B(n4), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15362_2_lut.init = 16'h2222;
    LUT4 i15361_2_lut (.A(n1105[5]), .B(n4), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15361_2_lut.init = 16'h2222;
    LUT4 i15360_2_lut (.A(n1105[4]), .B(n4), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15360_2_lut.init = 16'h2222;
    LUT4 i15359_2_lut (.A(n1105[3]), .B(n4), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15359_2_lut.init = 16'h2222;
    LUT4 i15358_2_lut (.A(n1105[2]), .B(n4), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15358_2_lut.init = 16'h2222;
    LUT4 i15357_2_lut (.A(n1105[1]), .B(n4), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15357_2_lut.init = 16'h2222;
    CCU2D add_1766_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26793), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_17.INIT0 = 16'hd222;
    defparam add_1766_17.INIT1 = 16'h0000;
    defparam add_1766_17.INJECT1_0 = "NO";
    defparam add_1766_17.INJECT1_1 = "NO";
    CCU2D add_1766_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26792), 
          .COUT(n26793), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_15.INIT0 = 16'hd222;
    defparam add_1766_15.INIT1 = 16'hd222;
    defparam add_1766_15.INJECT1_0 = "NO";
    defparam add_1766_15.INJECT1_1 = "NO";
    LUT4 i15111_2_lut (.A(n1105[0]), .B(n4), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15111_2_lut.init = 16'h2222;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14358), .PD(n16639), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1766_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26791), 
          .COUT(n26792), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_13.INIT0 = 16'hd222;
    defparam add_1766_13.INIT1 = 16'hd222;
    defparam add_1766_13.INJECT1_0 = "NO";
    defparam add_1766_13.INJECT1_1 = "NO";
    CCU2D add_1766_11 (.A0(\count[9] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26790), 
          .COUT(n26791), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_11.INIT0 = 16'hd222;
    defparam add_1766_11.INIT1 = 16'hd222;
    defparam add_1766_11.INJECT1_0 = "NO";
    defparam add_1766_11.INJECT1_1 = "NO";
    CCU2D add_1766_9 (.A0(\count[7] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26789), 
          .COUT(n26790), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_9.INIT0 = 16'hd222;
    defparam add_1766_9.INIT1 = 16'hd222;
    defparam add_1766_9.INJECT1_0 = "NO";
    defparam add_1766_9.INJECT1_1 = "NO";
    CCU2D add_1766_7 (.A0(\count[5] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26788), 
          .COUT(n26789), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1766_7.INIT0 = 16'hd222;
    defparam add_1766_7.INIT1 = 16'hd222;
    defparam add_1766_7.INJECT1_0 = "NO";
    defparam add_1766_7.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (n1168, n1180, n31964, GND_net, n30426, debug_c_c, 
            n31906, n33687, \register[2] , n14369, n1174, n27757, 
            n33685, n33686, rc_ch2_c, n29866) /* synthesis syn_module_defined=1 */ ;
    output n1168;
    output n1180;
    output n31964;
    input GND_net;
    output n30426;
    input debug_c_c;
    input n31906;
    input n33687;
    output [7:0]\register[2] ;
    input n14369;
    output n1174;
    input n27757;
    input n33685;
    input n33686;
    input rc_ch2_c;
    output n29866;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n32060, n29993, n27057;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    wire [7:0]n1096;
    
    wire n27056, n13395, n31994, n31967, n29219, n31969, n31995, 
        n22170, n27611, n31934, n31968, n27055, n27054, n27921, 
        n32066, n4, n32067, n4_adj_152;
    wire [15:0]n116;
    
    wire n16650;
    wire [7:0]n43;
    
    wire n29992, n29659, n22195, n31935, n6, n13472, n29925, n55, 
        n30251, n30184, n6_adj_153, n27867, n29926, n26801, n26800, 
        n26799, n26798, n26797, n26796, n26795, n26794;
    
    LUT4 i5_2_lut_rep_443 (.A(n1168), .B(n1180), .Z(n32060)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_443.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n1168), .B(n1180), .C(n31964), .Z(n29993)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    CCU2D sub_75_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27057), 
          .S0(n1096[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_9.INIT1 = 16'h0000;
    defparam sub_75_add_2_9.INJECT1_0 = "NO";
    defparam sub_75_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27056), 
          .COUT(n27057), .S0(n1096[5]), .S1(n1096[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_7.INJECT1_0 = "NO";
    defparam sub_75_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_377 (.A(count[9]), .B(n13395), .Z(n31994)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_377.init = 16'heeee;
    LUT4 i1_2_lut_rep_350_3_lut (.A(count[9]), .B(n13395), .C(count[8]), 
         .Z(n31967)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_350_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_352_4_lut (.A(count[9]), .B(n13395), .C(n29219), 
         .D(count[8]), .Z(n31969)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i2_3_lut_rep_352_4_lut.init = 16'hfeff;
    LUT4 i15567_2_lut_3_lut_4_lut (.A(count[9]), .B(n13395), .C(n31995), 
         .D(count[8]), .Z(n22170)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i15567_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_317_3_lut_4_lut (.A(count[9]), .B(n13395), .C(n27611), 
         .D(count[8]), .Z(n31934)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_317_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_378 (.A(count[0]), .B(n29219), .Z(n31995)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_378.init = 16'h8888;
    LUT4 i1_2_lut_rep_351_3_lut (.A(count[0]), .B(n29219), .C(count[8]), 
         .Z(n31968)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_351_3_lut.init = 16'h8080;
    CCU2D sub_75_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27055), 
          .COUT(n27056), .S0(n1096[3]), .S1(n1096[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_5.INJECT1_0 = "NO";
    defparam sub_75_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27054), 
          .COUT(n27055), .S0(n1096[1]), .S1(n1096[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_3.INJECT1_0 = "NO";
    defparam sub_75_add_2_3.INJECT1_1 = "NO";
    LUT4 i23114_2_lut_3_lut (.A(n1180), .B(n1168), .C(n27921), .Z(n30426)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i23114_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_449 (.A(count[6]), .B(count[7]), .Z(n32066)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_449.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_285 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_adj_285.init = 16'h8080;
    CCU2D sub_75_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27054), 
          .S1(n1096[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_1.INIT0 = 16'hF000;
    defparam sub_75_add_2_1.INIT1 = 16'h5555;
    defparam sub_75_add_2_1.INJECT1_0 = "NO";
    defparam sub_75_add_2_1.INJECT1_1 = "NO";
    LUT4 i3203_2_lut_rep_450 (.A(count[1]), .B(count[2]), .Z(n32067)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3203_2_lut_rep_450.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_286 (.A(count[1]), .B(count[2]), .C(count[3]), 
         .Z(n4_adj_152)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_286.init = 16'hf8f8;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31906), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31906), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31906), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31906), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31906), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31906), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31906), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31906), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33687), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33687), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3AX valid_48 (.D(n29992), .SP(n27757), .CK(debug_c_c), .Q(n1174));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(n1168), .B(n33685), .C(n29659), .D(n22195), .Z(n16650)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h0080;
    LUT4 i2_4_lut (.A(count[9]), .B(n27921), .C(n31968), .D(n1180), 
         .Z(n29659)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h00c8;
    LUT4 i23182_3_lut_3_lut_4_lut (.A(n27611), .B(n31967), .C(n22195), 
         .D(n31964), .Z(n29992)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23182_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i2_4_lut_adj_287 (.A(n31935), .B(n31969), .C(n31934), .D(n22170), 
         .Z(n27921)) /* synthesis lut_function=(A+!(B ((D)+!C))) */ ;
    defparam i2_4_lut_adj_287.init = 16'hbbfb;
    LUT4 i2_3_lut_4_lut (.A(n31968), .B(n22195), .C(n31994), .D(n31969), 
         .Z(n6)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_288 (.A(count[12]), .B(count[13]), .C(n13472), .D(n29925), 
         .Z(n13395)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_288.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[15]), .B(count[14]), .Z(n13472)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_289 (.A(count[11]), .B(count[10]), .Z(n29925)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_289.init = 16'heeee;
    LUT4 i2_4_lut_adj_290 (.A(count[4]), .B(n32066), .C(n4_adj_152), .D(count[5]), 
         .Z(n27611)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_290.init = 16'hc800;
    LUT4 i15592_4_lut (.A(count[9]), .B(n13395), .C(n55), .D(n30251), 
         .Z(n22195)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i15592_4_lut.init = 16'heeec;
    LUT4 i2_3_lut (.A(count[8]), .B(count[6]), .C(count[7]), .Z(n55)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i22841_4_lut (.A(count[5]), .B(count[3]), .C(count[4]), .D(n30184), 
         .Z(n30251)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i22841_4_lut.init = 16'ha080;
    LUT4 i22776_3_lut (.A(count[2]), .B(count[1]), .C(count[0]), .Z(n30184)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22776_3_lut.init = 16'hfefe;
    LUT4 i4_4_lut (.A(n32066), .B(count[1]), .C(count[3]), .D(n6_adj_153), 
         .Z(n29219)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h8000;
    LUT4 i1_3_lut (.A(count[2]), .B(count[5]), .C(count[4]), .Z(n6_adj_153)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_3_lut.init = 16'h8080;
    FD1P3AX prev_in_46 (.D(n1180), .SP(n33686), .CK(debug_c_c), .Q(n1168));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n33686), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1180));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_291 (.A(n31967), .B(n6), .C(n31995), .D(n27611), 
         .Z(n29866)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_291.init = 16'hc888;
    LUT4 i2_4_lut_adj_292 (.A(n29925), .B(n27867), .C(count[9]), .D(n4), 
         .Z(n29926)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i2_4_lut_adj_292.init = 16'hfefa;
    LUT4 i2_4_lut_adj_293 (.A(count[5]), .B(count[4]), .C(n32067), .D(count[3]), 
         .Z(n27867)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_293.init = 16'hfeee;
    CCU2D add_1762_17 (.A0(count[15]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26801), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_17.INIT0 = 16'hd222;
    defparam add_1762_17.INIT1 = 16'h0000;
    defparam add_1762_17.INJECT1_0 = "NO";
    defparam add_1762_17.INJECT1_1 = "NO";
    CCU2D add_1762_15 (.A0(count[13]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32060), .C1(GND_net), .D1(GND_net), .CIN(n26800), 
          .COUT(n26801), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_15.INIT0 = 16'hd222;
    defparam add_1762_15.INIT1 = 16'hd222;
    defparam add_1762_15.INJECT1_0 = "NO";
    defparam add_1762_15.INJECT1_1 = "NO";
    CCU2D add_1762_13 (.A0(count[11]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32060), .C1(GND_net), .D1(GND_net), .CIN(n26799), 
          .COUT(n26800), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_13.INIT0 = 16'hd222;
    defparam add_1762_13.INIT1 = 16'hd222;
    defparam add_1762_13.INJECT1_0 = "NO";
    defparam add_1762_13.INJECT1_1 = "NO";
    CCU2D add_1762_11 (.A0(count[9]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32060), .C1(GND_net), .D1(GND_net), .CIN(n26798), 
          .COUT(n26799), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_11.INIT0 = 16'hd222;
    defparam add_1762_11.INIT1 = 16'hd222;
    defparam add_1762_11.INJECT1_0 = "NO";
    defparam add_1762_11.INJECT1_1 = "NO";
    CCU2D add_1762_9 (.A0(count[7]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32060), .C1(GND_net), .D1(GND_net), .CIN(n26797), 
          .COUT(n26798), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_9.INIT0 = 16'hd222;
    defparam add_1762_9.INIT1 = 16'hd222;
    defparam add_1762_9.INJECT1_0 = "NO";
    defparam add_1762_9.INJECT1_1 = "NO";
    CCU2D add_1762_7 (.A0(count[5]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32060), .C1(GND_net), .D1(GND_net), .CIN(n26796), 
          .COUT(n26797), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_7.INIT0 = 16'hd222;
    defparam add_1762_7.INIT1 = 16'hd222;
    defparam add_1762_7.INJECT1_0 = "NO";
    defparam add_1762_7.INJECT1_1 = "NO";
    CCU2D add_1762_5 (.A0(count[3]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32060), .C1(GND_net), .D1(GND_net), .CIN(n26795), 
          .COUT(n26796), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_5.INIT0 = 16'hd222;
    defparam add_1762_5.INIT1 = 16'hd222;
    defparam add_1762_5.INJECT1_0 = "NO";
    defparam add_1762_5.INJECT1_1 = "NO";
    CCU2D add_1762_3 (.A0(count[1]), .B0(n32060), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32060), .C1(GND_net), .D1(GND_net), .CIN(n26794), 
          .COUT(n26795), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_3.INIT0 = 16'hd222;
    defparam add_1762_3.INIT1 = 16'hd222;
    defparam add_1762_3.INJECT1_0 = "NO";
    defparam add_1762_3.INJECT1_1 = "NO";
    CCU2D add_1762_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29993), .B1(n1180), .C1(count[0]), .D1(n1168), .COUT(n26794), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1762_1.INIT0 = 16'hF000;
    defparam add_1762_1.INIT1 = 16'ha565;
    defparam add_1762_1.INJECT1_0 = "NO";
    defparam add_1762_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14369), .PD(n16650), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i22710_4_lut_rep_347 (.A(n13472), .B(count[13]), .C(count[12]), 
         .D(n29926), .Z(n31964)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i22710_4_lut_rep_347.init = 16'heaaa;
    LUT4 i21_3_lut_rep_318_4_lut (.A(count[8]), .B(n31995), .C(n31994), 
         .D(n22195), .Z(n31935)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21_3_lut_rep_318_4_lut.init = 16'h00f8;
    LUT4 i15356_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15356_2_lut_4_lut.init = 16'h0400;
    LUT4 i15355_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15355_2_lut_4_lut.init = 16'h0400;
    LUT4 i15354_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15354_2_lut_4_lut.init = 16'h0400;
    LUT4 i15353_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15353_2_lut_4_lut.init = 16'h0400;
    LUT4 i15352_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15352_2_lut_4_lut.init = 16'h0400;
    LUT4 i15351_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15351_2_lut_4_lut.init = 16'h0400;
    LUT4 i15350_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15350_2_lut_4_lut.init = 16'h0400;
    LUT4 i15108_2_lut_4_lut (.A(n31994), .B(count[8]), .C(n29219), .D(n1096[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15108_2_lut_4_lut.init = 16'h0400;
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (GND_net, n1153, debug_c_c, n33686, n1165, n31948, 
            n30378, \register[1] , n14374, n33685, rc_ch1_c, n1159, 
            n27960, n29869) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n1153;
    input debug_c_c;
    input n33686;
    output n1165;
    output n31948;
    output n30378;
    output [7:0]\register[1] ;
    input n14374;
    input n33685;
    input rc_ch1_c;
    output n1159;
    input n27960;
    output n29869;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n29877, n6, n29879, n95;
    wire [7:0]n1087;
    
    wire n23;
    wire [7:0]n43;
    
    wire n27061, n27060, n27059, n27058, n31947, n22193, n32002, 
        n30200, n31980, n29930, n26809, n32082;
    wire [15:0]n116;
    
    wire n26808, n26807, n31979, n31927, n26806, n26805, n13384, 
        n31946, n27955, n4, n16653, n29929, n29657, n49_adj_151, 
        n30240, n26804, n30192, n26803, n13475, n29967, n26802, 
        n22176, n27892, n29968;
    
    LUT4 i1_4_lut (.A(count[4]), .B(n29877), .C(count[3]), .D(n6), .Z(n29879)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut.init = 16'hccc8;
    LUT4 i3261_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3261_2_lut.init = 16'h8888;
    LUT4 i3_4_lut (.A(count[3]), .B(count[4]), .C(count[2]), .D(n29877), 
         .Z(n95)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i15348_2_lut (.A(n1087[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15348_2_lut.init = 16'h8888;
    LUT4 i15347_2_lut (.A(n1087[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15347_2_lut.init = 16'h8888;
    LUT4 i15346_2_lut (.A(n1087[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15346_2_lut.init = 16'h8888;
    LUT4 i15345_2_lut (.A(n1087[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15345_2_lut.init = 16'h8888;
    LUT4 i15344_2_lut (.A(n1087[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15344_2_lut.init = 16'h8888;
    LUT4 i15343_2_lut (.A(n1087[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15343_2_lut.init = 16'h8888;
    CCU2D sub_74_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27061), 
          .S0(n1087[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_9.INIT1 = 16'h0000;
    defparam sub_74_add_2_9.INJECT1_0 = "NO";
    defparam sub_74_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27060), 
          .COUT(n27061), .S0(n1087[5]), .S1(n1087[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_7.INJECT1_0 = "NO";
    defparam sub_74_add_2_7.INJECT1_1 = "NO";
    FD1P3AX prev_in_46 (.D(n1165), .SP(n33686), .CK(debug_c_c), .Q(n1153));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D sub_74_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27059), 
          .COUT(n27060), .S0(n1087[3]), .S1(n1087[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_5.INJECT1_0 = "NO";
    defparam sub_74_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27058), 
          .COUT(n27059), .S0(n1087[1]), .S1(n1087[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_3.INJECT1_0 = "NO";
    defparam sub_74_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27058), 
          .S1(n1087[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_1.INIT0 = 16'hF000;
    defparam sub_74_add_2_1.INIT1 = 16'h5555;
    defparam sub_74_add_2_1.INJECT1_0 = "NO";
    defparam sub_74_add_2_1.INJECT1_1 = "NO";
    LUT4 i22792_3_lut_4_lut (.A(n31947), .B(n22193), .C(n32002), .D(n23), 
         .Z(n30200)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i22792_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23176_3_lut_3_lut_4_lut (.A(n29879), .B(n31980), .C(n22193), 
         .D(n31948), .Z(n29930)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23176_3_lut_3_lut_4_lut.init = 16'h000e;
    CCU2D add_1758_17 (.A0(count[15]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26809), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_17.INIT0 = 16'hd222;
    defparam add_1758_17.INIT1 = 16'h0000;
    defparam add_1758_17.INJECT1_0 = "NO";
    defparam add_1758_17.INJECT1_1 = "NO";
    CCU2D add_1758_15 (.A0(count[13]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32082), .C1(GND_net), .D1(GND_net), .CIN(n26808), 
          .COUT(n26809), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_15.INIT0 = 16'hd222;
    defparam add_1758_15.INIT1 = 16'hd222;
    defparam add_1758_15.INJECT1_0 = "NO";
    defparam add_1758_15.INJECT1_1 = "NO";
    CCU2D add_1758_13 (.A0(count[11]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32082), .C1(GND_net), .D1(GND_net), .CIN(n26807), 
          .COUT(n26808), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_13.INIT0 = 16'hd222;
    defparam add_1758_13.INIT1 = 16'hd222;
    defparam add_1758_13.INJECT1_0 = "NO";
    defparam add_1758_13.INJECT1_1 = "NO";
    LUT4 i21_3_lut_rep_310_4_lut (.A(count[8]), .B(n31979), .C(n32002), 
         .D(n22193), .Z(n31927)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21_3_lut_rep_310_4_lut.init = 16'h00f8;
    CCU2D add_1758_11 (.A0(count[9]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32082), .C1(GND_net), .D1(GND_net), .CIN(n26806), 
          .COUT(n26807), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_11.INIT0 = 16'hd222;
    defparam add_1758_11.INIT1 = 16'hd222;
    defparam add_1758_11.INJECT1_0 = "NO";
    defparam add_1758_11.INJECT1_1 = "NO";
    CCU2D add_1758_9 (.A0(count[7]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32082), .C1(GND_net), .D1(GND_net), .CIN(n26805), 
          .COUT(n26806), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_9.INIT0 = 16'hd222;
    defparam add_1758_9.INIT1 = 16'hd222;
    defparam add_1758_9.INJECT1_0 = "NO";
    defparam add_1758_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_385 (.A(count[9]), .B(n13384), .Z(n32002)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_385.init = 16'heeee;
    LUT4 i1_2_lut_rep_363_3_lut (.A(count[9]), .B(n13384), .C(count[8]), 
         .Z(n31980)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_363_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_329_3_lut_4_lut (.A(count[9]), .B(n13384), .C(n29879), 
         .D(count[8]), .Z(n31946)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_329_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23066_2_lut_3_lut (.A(n1165), .B(n1153), .C(n27955), .Z(n30378)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i23066_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), .Z(n29877)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_275 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_adj_275.init = 16'h8080;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i5_2_lut_rep_465 (.A(n1153), .B(n1165), .Z(n32082)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_465.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_276 (.A(n1153), .B(n1165), .C(n31948), .Z(n29929)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_adj_276.init = 16'hf4f4;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_277 (.A(n1153), .B(n33685), .C(n29657), .D(n22193), 
         .Z(n16653)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_277.init = 16'h0080;
    LUT4 i2_4_lut (.A(n31947), .B(n27955), .C(count[9]), .D(n1165), 
         .Z(n29657)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h00c8;
    LUT4 i15349_2_lut (.A(n1087[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15349_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_278 (.A(count[8]), .B(n32002), .C(count[1]), .D(n95), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_278.init = 16'h0222;
    LUT4 i15590_4_lut (.A(count[9]), .B(n13384), .C(n49_adj_151), .D(n30240), 
         .Z(n22193)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i15590_4_lut.init = 16'heeec;
    CCU2D add_1758_7 (.A0(count[5]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32082), .C1(GND_net), .D1(GND_net), .CIN(n26804), 
          .COUT(n26805), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_7.INIT0 = 16'hd222;
    defparam add_1758_7.INIT1 = 16'hd222;
    defparam add_1758_7.INJECT1_0 = "NO";
    defparam add_1758_7.INJECT1_1 = "NO";
    LUT4 i2_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n49_adj_151)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i22832_4_lut (.A(count[4]), .B(count[1]), .C(count[5]), .D(n30192), 
         .Z(n30240)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i22832_4_lut.init = 16'ha080;
    LUT4 i22784_3_lut (.A(count[0]), .B(count[2]), .C(count[3]), .Z(n30192)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22784_3_lut.init = 16'hfefe;
    CCU2D add_1758_5 (.A0(count[3]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32082), .C1(GND_net), .D1(GND_net), .CIN(n26803), 
          .COUT(n26804), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_5.INIT0 = 16'hd222;
    defparam add_1758_5.INIT1 = 16'hd222;
    defparam add_1758_5.INJECT1_0 = "NO";
    defparam add_1758_5.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_279 (.A(count[12]), .B(count[13]), .C(n13475), .D(n29967), 
         .Z(n13384)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_279.init = 16'hfffe;
    CCU2D add_1758_3 (.A0(count[1]), .B0(n32082), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32082), .C1(GND_net), .D1(GND_net), .CIN(n26802), 
          .COUT(n26803), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_3.INIT0 = 16'hd222;
    defparam add_1758_3.INIT1 = 16'hd222;
    defparam add_1758_3.INJECT1_0 = "NO";
    defparam add_1758_3.INJECT1_1 = "NO";
    CCU2D add_1758_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29929), .B1(n1165), .C1(count[0]), .D1(n1153), .COUT(n26802), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1758_1.INIT0 = 16'hF000;
    defparam add_1758_1.INIT1 = 16'ha565;
    defparam add_1758_1.INJECT1_0 = "NO";
    defparam add_1758_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(count[15]), .B(count[14]), .Z(n13475)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_280 (.A(count[10]), .B(count[11]), .Z(n29967)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_280.init = 16'heeee;
    LUT4 i2_4_lut_adj_281 (.A(n31927), .B(n23), .C(n31946), .D(n22176), 
         .Z(n27955)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_281.init = 16'heefe;
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n33686), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1165));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_362 (.A(n95), .B(count[1]), .C(count[0]), .Z(n31979)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_3_lut_rep_362.init = 16'h8080;
    LUT4 i15105_2_lut (.A(n1087[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15105_2_lut.init = 16'h8888;
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14374), .PD(n16653), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33686), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33686), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3AX valid_48 (.D(n29930), .SP(n27960), .CK(debug_c_c), .Q(n1159));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_330_4_lut (.A(n95), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n31947)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_330_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_282 (.A(n31980), .B(n30200), .C(n31979), .D(n29879), 
         .Z(n29869)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut_adj_282.init = 16'h3222;
    LUT4 i15573_2_lut_4_lut (.A(n95), .B(count[1]), .C(count[0]), .D(n31980), 
         .Z(n22176)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i15573_2_lut_4_lut.init = 16'hff80;
    LUT4 i2_4_lut_adj_283 (.A(n29967), .B(count[9]), .C(n27892), .D(n4), 
         .Z(n29968)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_283.init = 16'hfeee;
    LUT4 i2_4_lut_adj_284 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n27892)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_284.init = 16'hfeee;
    LUT4 i1_4_lut_rep_331 (.A(n13475), .B(count[13]), .C(count[12]), .D(n29968), 
         .Z(n31948)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_331.init = 16'heaaa;
    
endmodule
//
// Verilog Description of module SabertoothSerialPeripheral
//

module SabertoothSerialPeripheral (debug_c_c, n13557, n282, n31991, 
            \databus[6] , \databus[5] , \databus[4] , \databus[3] , 
            \databus[2] , \databus[1] , \databus[0] , \register[0] , 
            n22326, \read_size[0] , n31922, \select[2] , n9366, rw, 
            n32075, n31940, \register_addr[0] , \reset_count[14] , n22296, 
            n5, n5_adj_44, n5_adj_45, n5_adj_46, n5_adj_47, n5_adj_48, 
            n5_adj_49, n32088, n89, n5_adj_50, \state[0] , GND_net, 
            n12, n31907, n7, n31908, n18379, n5497, n18374, n5495, 
            n5494, n5493, n32016, n29, \state[1] , n7648, n92, 
            n25, n94, n27, n93, n26, n91, n28, n90, n30, \reset_count[6] , 
            \reset_count[5] , \reset_count[4] , n47, \reset_count[8] , 
            \reset_count[7] , n29946, \state[3] , \state[2] , n31515, 
            \reset_count[11] , n21480, n27577, n29900, n14519, n31957, 
            motor_pwm_l_c, n8343, n2954, n30355, select_clk, n107) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n13557;
    input n282;
    input n31991;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    input \databus[0] ;
    output [7:0]\register[0] ;
    input n22326;
    output \read_size[0] ;
    input n31922;
    input \select[2] ;
    input n9366;
    input rw;
    output n32075;
    input n31940;
    input \register_addr[0] ;
    input \reset_count[14] ;
    input n22296;
    output n5;
    output n5_adj_44;
    output n5_adj_45;
    output n5_adj_46;
    output n5_adj_47;
    output n5_adj_48;
    output n5_adj_49;
    input n32088;
    output n89;
    output n5_adj_50;
    output \state[0] ;
    input GND_net;
    input n12;
    input n31907;
    output n7;
    input n31908;
    input n18379;
    input n5497;
    input n18374;
    input n5495;
    input n5494;
    input n5493;
    input n32016;
    output n29;
    output \state[1] ;
    input n7648;
    output n92;
    output n25;
    output n94;
    output n27;
    output n93;
    output n26;
    output n91;
    output n28;
    output n90;
    output n30;
    input \reset_count[6] ;
    input \reset_count[5] ;
    input \reset_count[4] ;
    output n47;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29946;
    output \state[3] ;
    output \state[2] ;
    output n31515;
    input \reset_count[11] ;
    input n21480;
    input n27577;
    output n29900;
    input n14519;
    input n31957;
    output motor_pwm_l_c;
    output n8343;
    input n2954;
    output n30355;
    output select_clk;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n31916;
    wire [7:0]\register[0]_c ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n31912, n14675, prev_select;
    wire [7:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(92[12:22])
    wire [7:0]n1;
    
    wire n30032, n9277, n32015, n27635, n9274;
    wire [7:0]n6182;
    
    FD1P3AX register_0__i16 (.D(n282), .SP(n13557), .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n31916), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n31916), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n31916), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n31916), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n31916), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n31916), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n31916), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n282), .SP(n22326), .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n31912), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[0]_c [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n31912), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[0]_c [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n31912), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[0]_c [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n31912), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[0]_c [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n31912), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[0]_c [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n31912), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[0]_c [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i2.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n31922), .SP(n14675), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n31912), .PD(n31991), 
            .CK(debug_c_c), .Q(\register[0]_c [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam prev_select_138.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n1[0]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i23078_2_lut_rep_295_4_lut (.A(rw), .B(n32075), .C(n31940), .D(\register_addr[0] ), 
         .Z(n31912)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i23078_2_lut_rep_295_4_lut.init = 16'h0004;
    LUT4 i4538_2_lut_rep_299_4_lut (.A(rw), .B(n32075), .C(n31940), .D(\register_addr[0] ), 
         .Z(n31916)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i4538_2_lut_rep_299_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_458 (.A(\select[2] ), .B(prev_select), .Z(n32075)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_rep_458.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\select[2] ), .B(prev_select), .C(\reset_count[14] ), 
         .D(n22296), .Z(n14675)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4247_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[7]), 
         .Z(n5)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4247_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4248_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[6]), 
         .Z(n5_adj_44)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4248_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4249_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[5]), 
         .Z(n5_adj_45)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4249_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4250_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[4]), 
         .Z(n5_adj_46)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4250_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4251_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[3]), 
         .Z(n5_adj_47)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4251_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4254_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[0]), 
         .Z(n5_adj_48)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4254_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4253_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[1]), 
         .Z(n5_adj_49)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4253_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 i15341_4_lut_4_lut (.A(\register[1] [7]), .B(n32088), .C(n30032), 
         .D(n9277), .Z(n89)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i15341_4_lut_4_lut.init = 16'hffde;
    LUT4 i1_4_lut_4_lut (.A(\register[1] [7]), .B(n32088), .C(\register[1] [1]), 
         .D(n32015), .Z(n9277)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i1_4_lut_4_lut.init = 16'h2000;
    LUT4 Select_4252_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[2]), 
         .Z(n5_adj_50)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4252_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_4_lut_adj_274 (.A(\register[0] [7]), .B(n32088), .C(\register[0]_c [1]), 
         .D(n27635), .Z(n9274)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i1_4_lut_4_lut_adj_274.init = 16'h2000;
    LUT4 mux_1899_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n6182[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1899_Mux_6_i1_3_lut (.A(\register[0]_c [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n6182[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1899_Mux_5_i1_3_lut (.A(\register[0]_c [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n6182[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1899_Mux_4_i1_3_lut (.A(\register[0]_c [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n6182[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1899_Mux_3_i1_3_lut (.A(\register[0]_c [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n6182[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1899_Mux_2_i1_3_lut (.A(\register[0]_c [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n6182[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1899_Mux_1_i1_3_lut (.A(\register[0]_c [1]), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n6182[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_1_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i7 (.D(n6182[7]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6182[6]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6182[5]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6182[4]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6182[3]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n6182[2]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n6182[1]), .SP(n14675), .CD(n9366), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=534, LSE_RLINE=542 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1899_Mux_0_i1_3_lut (.A(\register[0]_c [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n1[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1899_Mux_0_i1_3_lut.init = 16'hcaca;
    SabertoothSerial sserial (.\state[0] (\state[0] ), .debug_c_c(debug_c_c), 
            .GND_net(GND_net), .n12(n12), .\register[0][1] (\register[0]_c [1]), 
            .n27635(n27635), .\register[0][7] (\register[0] [7]), .\register[0][4] (\register[0]_c [4]), 
            .\register[0][6] (\register[0]_c [6]), .\register[0][5] (\register[0]_c [5]), 
            .\register[1][4] (\register[1] [4]), .\register[1][6] (\register[1] [6]), 
            .\register[1][5] (\register[1] [5]), .n30032(n30032), .\register[0][2] (\register[0]_c [2]), 
            .\register[0][3] (\register[0]_c [3]), .\register[1][2] (\register[1] [2]), 
            .\register[1][1] (\register[1] [1]), .\register[1][3] (\register[1] [3]), 
            .n31907(n31907), .n7(n7), .n32088(n32088), .n32015(n32015), 
            .\register[1][7] (\register[1] [7]), .n31908(n31908), .n18379(n18379), 
            .n5497(n5497), .n18374(n18374), .n5495(n5495), .n5494(n5494), 
            .n5493(n5493), .n32016(n32016), .n9274(n9274), .n29(n29), 
            .\state[1] (\state[1] ), .n7648(n7648), .n9277(n9277), .n92(n92), 
            .n25(n25), .n94(n94), .n27(n27), .n93(n93), .n26(n26), 
            .n91(n91), .n28(n28), .n90(n90), .n30(n30), .n31991(n31991), 
            .\reset_count[6] (\reset_count[6] ), .\reset_count[5] (\reset_count[5] ), 
            .\reset_count[4] (\reset_count[4] ), .n47(n47), .\reset_count[8] (\reset_count[8] ), 
            .\reset_count[7] (\reset_count[7] ), .n29946(n29946), .\state[3] (\state[3] ), 
            .\state[2] (\state[2] ), .n31515(n31515), .\reset_count[11] (\reset_count[11] ), 
            .n21480(n21480), .n27577(n27577), .n29900(n29900), .n14519(n14519), 
            .n31957(n31957), .motor_pwm_l_c(motor_pwm_l_c), .n22296(n22296), 
            .\reset_count[14] (\reset_count[14] ), .n8343(n8343), .n2954(n2954), 
            .n30355(n30355), .select_clk(select_clk), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(142[19] 147[34])
    
endmodule
//
// Verilog Description of module SabertoothSerial
//

module SabertoothSerial (\state[0] , debug_c_c, GND_net, n12, \register[0][1] , 
            n27635, \register[0][7] , \register[0][4] , \register[0][6] , 
            \register[0][5] , \register[1][4] , \register[1][6] , \register[1][5] , 
            n30032, \register[0][2] , \register[0][3] , \register[1][2] , 
            \register[1][1] , \register[1][3] , n31907, n7, n32088, 
            n32015, \register[1][7] , n31908, n18379, n5497, n18374, 
            n5495, n5494, n5493, n32016, n9274, n29, \state[1] , 
            n7648, n9277, n92, n25, n94, n27, n93, n26, n91, 
            n28, n90, n30, n31991, \reset_count[6] , \reset_count[5] , 
            \reset_count[4] , n47, \reset_count[8] , \reset_count[7] , 
            n29946, \state[3] , \state[2] , n31515, \reset_count[11] , 
            n21480, n27577, n29900, n14519, n31957, motor_pwm_l_c, 
            n22296, \reset_count[14] , n8343, n2954, n30355, select_clk, 
            n107) /* synthesis syn_module_defined=1 */ ;
    output \state[0] ;
    input debug_c_c;
    input GND_net;
    input n12;
    input \register[0][1] ;
    output n27635;
    input \register[0][7] ;
    input \register[0][4] ;
    input \register[0][6] ;
    input \register[0][5] ;
    input \register[1][4] ;
    input \register[1][6] ;
    input \register[1][5] ;
    output n30032;
    input \register[0][2] ;
    input \register[0][3] ;
    input \register[1][2] ;
    input \register[1][1] ;
    input \register[1][3] ;
    input n31907;
    output n7;
    input n32088;
    output n32015;
    input \register[1][7] ;
    input n31908;
    input n18379;
    input n5497;
    input n18374;
    input n5495;
    input n5494;
    input n5493;
    input n32016;
    input n9274;
    output n29;
    output \state[1] ;
    input n7648;
    input n9277;
    output n92;
    output n25;
    output n94;
    output n27;
    output n93;
    output n26;
    output n91;
    output n28;
    output n90;
    output n30;
    input n31991;
    input \reset_count[6] ;
    input \reset_count[5] ;
    input \reset_count[4] ;
    output n47;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29946;
    output \state[3] ;
    output \state[2] ;
    output n31515;
    input \reset_count[11] ;
    input n21480;
    input n27577;
    output n29900;
    input n14519;
    input n31957;
    output motor_pwm_l_c;
    input n22296;
    input \reset_count[14] ;
    output n8343;
    input n2954;
    output n30355;
    output select_clk;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n40, n24, n32013, n12514, n32014, n32054, n11805, n31988, 
        n11908, n32055, n31989;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(16[12:19])
    
    wire n31901, n20, n31956, n12516, n31954, n29761, n1150, n1, 
        n29590, n6, n28668, n10146, n6_adj_142, n8, n12_adj_143, 
        n11778;
    
    FD1S3IX state__i0 (.D(n12), .CK(debug_c_c), .CD(GND_net), .Q(\state[0] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n40), .B(\register[0][1] ), .C(n27635), .D(\register[0][7] ), 
         .Z(n24)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;
    defparam i1_4_lut.init = 16'h5111;
    LUT4 i5884_2_lut_3_lut_4_lut (.A(\register[0][4] ), .B(n32013), .C(\register[0][6] ), 
         .D(\register[0][5] ), .Z(n12514)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5884_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i22630_2_lut_3_lut_4_lut (.A(\register[1][4] ), .B(n32014), .C(\register[1][6] ), 
         .D(\register[1][5] ), .Z(n30032)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22630_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i5164_2_lut_rep_437 (.A(\register[0][2] ), .B(\register[0][1] ), 
         .Z(n32054)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5164_2_lut_rep_437.init = 16'h8888;
    LUT4 i5168_2_lut_rep_396_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n32013)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5168_2_lut_rep_396_3_lut.init = 16'h8080;
    LUT4 i5179_2_lut_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n11805)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i5179_2_lut_3_lut.init = 16'h7878;
    LUT4 i5866_2_lut_rep_371_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n31988)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5866_2_lut_rep_371_3_lut_4_lut.init = 16'h8000;
    LUT4 i5282_2_lut_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n11908)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5282_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4390_2_lut_rep_438 (.A(\register[1][2] ), .B(\register[1][1] ), 
         .Z(n32055)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4390_2_lut_rep_438.init = 16'h8888;
    LUT4 i5736_2_lut_rep_372_3_lut_4_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][4] ), .D(\register[1][3] ), .Z(n31989)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5736_2_lut_rep_372_3_lut_4_lut.init = 16'h8000;
    LUT4 i4622_2_lut_rep_397_3_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][3] ), .Z(n32014)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i4622_2_lut_rep_397_3_lut.init = 16'h8080;
    FD1P3AX tx_data_i0_i0 (.D(n31901), .SP(n31907), .CK(debug_c_c), .Q(tx_data[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    LUT4 n20_bdd_4_lut (.A(n20), .B(n24), .C(n7), .D(n32088), .Z(n31901)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n20_bdd_4_lut.init = 16'h00ca;
    LUT4 i5868_2_lut_rep_339_3_lut_4_lut (.A(\register[0][3] ), .B(n32054), 
         .C(\register[0][5] ), .D(\register[0][4] ), .Z(n31956)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5868_2_lut_rep_339_3_lut_4_lut.init = 16'h8000;
    LUT4 i5886_2_lut_3_lut_4_lut (.A(\register[0][3] ), .B(n32054), .C(\register[0][5] ), 
         .D(\register[0][4] ), .Z(n12516)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5886_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i5850_2_lut_rep_337_3_lut_4_lut (.A(\register[1][3] ), .B(n32055), 
         .C(\register[1][5] ), .D(\register[1][4] ), .Z(n31954)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5850_2_lut_rep_337_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_398 (.A(\register[1][6] ), .B(n29761), .Z(n32015)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_398.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(\register[1][6] ), .B(n29761), .C(\register[1][7] ), 
         .D(\register[1][1] ), .Z(n20)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h80ff;
    FD1P3IX send_31 (.D(n1), .SP(n31908), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1150));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam send_31.GSR = "ENABLED";
    PFUMX i30 (.BLUT(n29590), .ALUT(n6), .C0(n7), .Z(n28668));
    LUT4 i3909_1_lut (.A(\state[0] ), .Z(n1)) /* synthesis lut_function=(!(A)) */ ;
    defparam i3909_1_lut.init = 16'h5555;
    LUT4 i14735_3_lut_4_lut (.A(\register[0][5] ), .B(n31988), .C(n32088), 
         .D(\register[0][6] ), .Z(n10146)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i14735_3_lut_4_lut.init = 16'hf8f0;
    FD1P3AX tx_data_i0_i1 (.D(n18379), .SP(n31907), .CK(debug_c_c), .Q(tx_data[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i2 (.D(n5497), .SP(n31907), .CK(debug_c_c), .Q(tx_data[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n18374), .SP(n31907), .CK(debug_c_c), .Q(tx_data[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n5495), .SP(n31907), .CK(debug_c_c), .Q(tx_data[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i5 (.D(n5494), .SP(n31907), .CK(debug_c_c), .Q(tx_data[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i6 (.D(n5493), .SP(n31907), .CK(debug_c_c), .Q(tx_data[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i7 (.D(n28668), .SP(n31907), .CK(debug_c_c), .Q(tx_data[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_266 (.A(n32016), .B(n40), .C(n9274), .D(n10146), 
         .Z(n29)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_266.init = 16'h3132;
    LUT4 equal_16_i5_2_lut (.A(\state[0] ), .B(\state[1] ), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(46[7:11])
    defparam equal_16_i5_2_lut.init = 16'hbbbb;
    LUT4 i40_2_lut (.A(\state[0] ), .B(\state[1] ), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i40_2_lut.init = 16'heeee;
    LUT4 i4_4_lut (.A(\register[0][4] ), .B(\register[0][2] ), .C(\register[0][3] ), 
         .D(n6_adj_142), .Z(n27635)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(\register[0][5] ), .B(\register[0][6] ), .Z(n6_adj_142)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i3_4_lut (.A(\register[1][4] ), .B(\register[1][3] ), .C(\register[1][5] ), 
         .D(\register[1][2] ), .Z(n29761)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    FD1P3IX state__i1 (.D(n7648), .SP(n31908), .CD(GND_net), .CK(debug_c_c), 
            .Q(\state[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_267 (.A(n32088), .B(\register[1][7] ), .C(n30032), 
         .D(n8), .Z(n29590)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_267.init = 16'hffbf;
    LUT4 i1_2_lut_adj_268 (.A(\register[1][1] ), .B(n29761), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_268.init = 16'h8888;
    LUT4 i6_4_lut (.A(n31956), .B(n12_adj_143), .C(\register[0][7] ), 
         .D(\state[1] ), .Z(n6)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i6_4_lut.init = 16'h0080;
    LUT4 i5_4_lut (.A(\register[0][6] ), .B(\state[0] ), .C(n9274), .D(n32088), 
         .Z(n12_adj_143)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i5_4_lut.init = 16'h0002;
    LUT4 i15338_4_lut (.A(\register[1][4] ), .B(n9277), .C(n32088), .D(n32014), 
         .Z(n92)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15338_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_269 (.A(n11908), .B(n40), .C(n9274), .D(n32088), 
         .Z(n25)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_269.init = 16'h3032;
    LUT4 i15336_4_lut (.A(\register[1][2] ), .B(n9277), .C(n32088), .D(\register[1][1] ), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15336_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_270 (.A(n11778), .B(n40), .C(n9274), .D(n32088), 
         .Z(n27)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_270.init = 16'h3032;
    LUT4 i5152_2_lut (.A(\register[0][2] ), .B(\register[0][1] ), .Z(n11778)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5152_2_lut.init = 16'h6666;
    LUT4 i15337_4_lut (.A(\register[1][3] ), .B(n9277), .C(n32088), .D(n32055), 
         .Z(n93)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15337_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_271 (.A(n11805), .B(n40), .C(n9274), .D(n32088), 
         .Z(n26)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_271.init = 16'h3032;
    LUT4 i15339_4_lut (.A(\register[1][5] ), .B(n9277), .C(n32088), .D(n31989), 
         .Z(n91)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15339_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_272 (.A(n12516), .B(n40), .C(n9274), .D(n32088), 
         .Z(n28)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_272.init = 16'h3032;
    LUT4 i15340_4_lut (.A(\register[1][6] ), .B(n9277), .C(n32088), .D(n31954), 
         .Z(n90)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15340_4_lut.init = 16'hcdce;
    LUT4 i1_4_lut_adj_273 (.A(n12514), .B(n40), .C(n9274), .D(n32088), 
         .Z(n30)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_4_lut_adj_273.init = 16'h3032;
    \UARTTransmitter(baud_div=1250)  sender (.n31991(n31991), .\reset_count[6] (\reset_count[6] ), 
            .\reset_count[5] (\reset_count[5] ), .\reset_count[4] (\reset_count[4] ), 
            .n47(n47), .\reset_count[8] (\reset_count[8] ), .\reset_count[7] (\reset_count[7] ), 
            .n29946(n29946), .\state[3] (\state[3] ), .\state[2] (\state[2] ), 
            .n1150(n1150), .n31515(n31515), .\reset_count[11] (\reset_count[11] ), 
            .n21480(n21480), .n27577(n27577), .n29900(n29900), .tx_data({tx_data}), 
            .n14519(n14519), .n31957(n31957), .motor_pwm_l_c(motor_pwm_l_c), 
            .n22296(n22296), .\reset_count[14] (\reset_count[14] ), .GND_net(GND_net), 
            .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(63[26] 67[47])
    \ClockDividerP(factor=12000)  baud_gen (.GND_net(GND_net), .n8343(n8343), 
            .debug_c_c(debug_c_c), .n2954(n2954), .n30355(n30355), .select_clk(select_clk), 
            .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(21[25] 23[48])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=1250) 
//

module \UARTTransmitter(baud_div=1250)  (n31991, \reset_count[6] , \reset_count[5] , 
            \reset_count[4] , n47, \reset_count[8] , \reset_count[7] , 
            n29946, \state[3] , \state[2] , n1150, n31515, \reset_count[11] , 
            n21480, n27577, n29900, tx_data, n14519, n31957, motor_pwm_l_c, 
            n22296, \reset_count[14] , GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input n31991;
    input \reset_count[6] ;
    input \reset_count[5] ;
    input \reset_count[4] ;
    output n47;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29946;
    output \state[3] ;
    output \state[2] ;
    input n1150;
    output n31515;
    input \reset_count[11] ;
    input n21480;
    input n27577;
    output n29900;
    input [7:0]tx_data;
    input n14519;
    input n31957;
    output motor_pwm_l_c;
    input n22296;
    input \reset_count[14] ;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n31079, n2773, n28780, n31077, n31076, n31078;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9281, n2, n30298, n7, n10, n29849, n104, n29850, n30296, 
        n30297, n10_adj_141, n21535;
    
    FD1S3IX state__i0 (.D(n31079), .CK(bclk), .CD(n31991), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(\reset_count[6] ), .B(\reset_count[5] ), .C(\reset_count[4] ), 
         .Z(n47)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i1_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut (.A(\reset_count[8] ), .B(\reset_count[7] ), .Z(n29946)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut (.A(n31991), .B(\state[3] ), .C(\state[2] ), .D(n2773), 
         .Z(n28780)) /* synthesis lut_function=(!(A+(B (C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h1404;
    LUT4 n1150_bdd_4_lut (.A(n1150), .B(state[1]), .C(\state[3] ), .D(state[0]), 
         .Z(n31515)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam n1150_bdd_4_lut.init = 16'h8001;
    LUT4 state_1__bdd_2_lut (.A(state[0]), .B(\state[3] ), .Z(n31077)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 state_0__bdd_4_lut (.A(state[0]), .B(state[1]), .C(\state[3] ), 
         .D(\state[2] ), .Z(n31076)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam state_0__bdd_4_lut.init = 16'h0f7e;
    LUT4 i1_4_lut_adj_264 (.A(\reset_count[11] ), .B(n21480), .C(\reset_count[8] ), 
         .D(n27577), .Z(n29900)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_264.init = 16'h8880;
    LUT4 state_1__bdd_4_lut_23720 (.A(state[1]), .B(state[0]), .C(n1150), 
         .D(\state[3] ), .Z(n31078)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;
    defparam state_1__bdd_4_lut_23720.init = 16'hb332;
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9281), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n30298), .C(\state[2] ), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15392_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15392_4_lut.init = 16'hfcee;
    FD1P3AX state__i3 (.D(n28780), .SP(n14519), .CK(bclk), .Q(\state[3] )) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(n31991), .B(\state[2] ), .C(\state[3] ), .D(n2773), 
         .Z(n29849)) /* synthesis lut_function=(!(A+(B (C+(D))+!B !(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1104;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(\state[3] ), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;
    LUT4 i1_3_lut_adj_265 (.A(state[1]), .B(n31957), .C(state[0]), .Z(n29850)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut_adj_265.init = 16'h4848;
    FD1P3AX state__i2 (.D(n29849), .SP(n14519), .CK(bclk), .Q(\state[2] )) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n29850), .SP(n14519), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3JX tx_35 (.D(n104), .SP(n31076), .PD(n31991), .CK(bclk), .Q(motor_pwm_l_c)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    PFUMX i22888 (.BLUT(n30296), .ALUT(n30297), .C0(state[1]), .Z(n30298));
    LUT4 i932_2_lut (.A(state[0]), .B(state[1]), .Z(n2773)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i932_2_lut.init = 16'h8888;
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9281), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9281), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9281), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9281), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9281), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9281), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9281), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i5_3_lut (.A(n22296), .B(n10_adj_141), .C(state[1]), .Z(n9281)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i5_3_lut.init = 16'h0808;
    PFUMX i23334 (.BLUT(n31078), .ALUT(n31077), .C0(\state[2] ), .Z(n31079));
    LUT4 i4_4_lut (.A(n21535), .B(\state[2] ), .C(n1150), .D(\reset_count[14] ), 
         .Z(n10_adj_141)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4_4_lut.init = 16'h1000;
    LUT4 i14941_2_lut (.A(\state[3] ), .B(state[0]), .Z(n21535)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14941_2_lut.init = 16'heeee;
    LUT4 i22886_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n30296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22886_3_lut.init = 16'hcaca;
    LUT4 i22887_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n30297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22887_3_lut.init = 16'hcaca;
    \ClockDividerP(factor=1250)  baud_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .bclk(bclk)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=1250) 
//

module \ClockDividerP(factor=1250)  (GND_net, debug_c_c, bclk) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    output bclk;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    
    wire n28110;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n8, n16541, n39, n52, n48, n40, n31, n50, n44, n32, 
        n42, n46, n36, n27427;
    wire [31:0]n102;
    
    wire n27426, n27425, n27424, n27423, n27422, n27421, n27420, 
        n27419, n27418, n27219, n8378, n27417, n27218, n27217, 
        n27416, n27216, n27215, n27415, n27214, n27213, n27414, 
        n27212, n27211, n27413, n27210, n27209, n27412, n27208, 
        n27207, n27206, n27205;
    
    LUT4 i23128_4_lut (.A(n28110), .B(count[5]), .C(n8), .D(count[0]), 
         .Z(n16541)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23128_4_lut.init = 16'h4000;
    LUT4 i26_4_lut (.A(n39), .B(n52), .C(n48), .D(n40), .Z(n28110)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i3_3_lut (.A(count[10]), .B(count[6]), .C(count[7]), .Z(n8)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3_3_lut.init = 16'h8080;
    LUT4 i12_2_lut (.A(count[30]), .B(count[13]), .Z(n39)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i12_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(n31), .B(n50), .C(n44), .D(n32), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(count[27]), .B(n42), .C(count[23]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(count[22]), .B(count[18]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i4_2_lut (.A(count[28]), .B(count[9]), .Z(n31)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(count[19]), .B(n46), .C(n36), .D(count[25]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(count[4]), .B(count[11]), .C(count[8]), .D(count[14]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[12]), .B(count[1]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[20]), .B(count[2]), .C(count[24]), .D(count[29]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(count[26]), .B(count[3]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i15_4_lut (.A(count[16]), .B(count[15]), .C(count[31]), .D(count[21]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_4_lut.init = 16'hfffe;
    CCU2D count_2643_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27427), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_33.INIT1 = 16'h0000;
    defparam count_2643_add_4_33.INJECT1_0 = "NO";
    defparam count_2643_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27426), .COUT(n27427), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_31.INJECT1_0 = "NO";
    defparam count_2643_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27425), .COUT(n27426), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_29.INJECT1_0 = "NO";
    defparam count_2643_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27424), .COUT(n27425), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_27.INJECT1_0 = "NO";
    defparam count_2643_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27423), .COUT(n27424), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_25.INJECT1_0 = "NO";
    defparam count_2643_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27422), .COUT(n27423), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_23.INJECT1_0 = "NO";
    defparam count_2643_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27421), .COUT(n27422), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_21.INJECT1_0 = "NO";
    defparam count_2643_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27420), .COUT(n27421), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_19.INJECT1_0 = "NO";
    defparam count_2643_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27419), .COUT(n27420), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_17.INJECT1_0 = "NO";
    defparam count_2643_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27418), .COUT(n27419), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_15.INJECT1_0 = "NO";
    defparam count_2643_add_4_15.INJECT1_1 = "NO";
    CCU2D add_20101_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27219), 
          .S1(n8378));
    defparam add_20101_32.INIT0 = 16'h5555;
    defparam add_20101_32.INIT1 = 16'h0000;
    defparam add_20101_32.INJECT1_0 = "NO";
    defparam add_20101_32.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27417), .COUT(n27418), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_13.INJECT1_0 = "NO";
    defparam count_2643_add_4_13.INJECT1_1 = "NO";
    CCU2D add_20101_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27218), .COUT(n27219));
    defparam add_20101_30.INIT0 = 16'h5555;
    defparam add_20101_30.INIT1 = 16'h5555;
    defparam add_20101_30.INJECT1_0 = "NO";
    defparam add_20101_30.INJECT1_1 = "NO";
    CCU2D add_20101_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27217), .COUT(n27218));
    defparam add_20101_28.INIT0 = 16'h5555;
    defparam add_20101_28.INIT1 = 16'h5555;
    defparam add_20101_28.INJECT1_0 = "NO";
    defparam add_20101_28.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27416), .COUT(n27417), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_11.INJECT1_0 = "NO";
    defparam count_2643_add_4_11.INJECT1_1 = "NO";
    CCU2D add_20101_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27216), .COUT(n27217));
    defparam add_20101_26.INIT0 = 16'h5555;
    defparam add_20101_26.INIT1 = 16'h5555;
    defparam add_20101_26.INJECT1_0 = "NO";
    defparam add_20101_26.INJECT1_1 = "NO";
    CCU2D add_20101_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27215), .COUT(n27216));
    defparam add_20101_24.INIT0 = 16'h5555;
    defparam add_20101_24.INIT1 = 16'h5555;
    defparam add_20101_24.INJECT1_0 = "NO";
    defparam add_20101_24.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27415), .COUT(n27416), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_9.INJECT1_0 = "NO";
    defparam count_2643_add_4_9.INJECT1_1 = "NO";
    CCU2D add_20101_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27214), .COUT(n27215));
    defparam add_20101_22.INIT0 = 16'h5555;
    defparam add_20101_22.INIT1 = 16'h5555;
    defparam add_20101_22.INJECT1_0 = "NO";
    defparam add_20101_22.INJECT1_1 = "NO";
    CCU2D add_20101_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27213), .COUT(n27214));
    defparam add_20101_20.INIT0 = 16'h5555;
    defparam add_20101_20.INIT1 = 16'h5555;
    defparam add_20101_20.INJECT1_0 = "NO";
    defparam add_20101_20.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27414), .COUT(n27415), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_7.INJECT1_0 = "NO";
    defparam count_2643_add_4_7.INJECT1_1 = "NO";
    CCU2D add_20101_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27212), .COUT(n27213));
    defparam add_20101_18.INIT0 = 16'h5555;
    defparam add_20101_18.INIT1 = 16'h5555;
    defparam add_20101_18.INJECT1_0 = "NO";
    defparam add_20101_18.INJECT1_1 = "NO";
    CCU2D add_20101_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27211), .COUT(n27212));
    defparam add_20101_16.INIT0 = 16'h5555;
    defparam add_20101_16.INIT1 = 16'h5555;
    defparam add_20101_16.INJECT1_0 = "NO";
    defparam add_20101_16.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27413), .COUT(n27414), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_5.INJECT1_0 = "NO";
    defparam count_2643_add_4_5.INJECT1_1 = "NO";
    CCU2D add_20101_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27210), .COUT(n27211));
    defparam add_20101_14.INIT0 = 16'h5555;
    defparam add_20101_14.INIT1 = 16'h5555;
    defparam add_20101_14.INJECT1_0 = "NO";
    defparam add_20101_14.INJECT1_1 = "NO";
    CCU2D add_20101_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27209), .COUT(n27210));
    defparam add_20101_12.INIT0 = 16'h5555;
    defparam add_20101_12.INIT1 = 16'h5555;
    defparam add_20101_12.INJECT1_0 = "NO";
    defparam add_20101_12.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27412), .COUT(n27413), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2643_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2643_add_4_3.INJECT1_0 = "NO";
    defparam count_2643_add_4_3.INJECT1_1 = "NO";
    CCU2D add_20101_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27208), .COUT(n27209));
    defparam add_20101_10.INIT0 = 16'h5aaa;
    defparam add_20101_10.INIT1 = 16'h5555;
    defparam add_20101_10.INJECT1_0 = "NO";
    defparam add_20101_10.INJECT1_1 = "NO";
    CCU2D add_20101_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27207), 
          .COUT(n27208));
    defparam add_20101_8.INIT0 = 16'h5555;
    defparam add_20101_8.INIT1 = 16'h5555;
    defparam add_20101_8.INJECT1_0 = "NO";
    defparam add_20101_8.INJECT1_1 = "NO";
    CCU2D add_20101_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27206), 
          .COUT(n27207));
    defparam add_20101_6.INIT0 = 16'h5aaa;
    defparam add_20101_6.INIT1 = 16'h5aaa;
    defparam add_20101_6.INJECT1_0 = "NO";
    defparam add_20101_6.INJECT1_1 = "NO";
    CCU2D count_2643_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27412), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643_add_4_1.INIT0 = 16'hF000;
    defparam count_2643_add_4_1.INIT1 = 16'h0555;
    defparam count_2643_add_4_1.INJECT1_0 = "NO";
    defparam count_2643_add_4_1.INJECT1_1 = "NO";
    CCU2D add_20101_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27205), 
          .COUT(n27206));
    defparam add_20101_4.INIT0 = 16'h5555;
    defparam add_20101_4.INIT1 = 16'h5aaa;
    defparam add_20101_4.INJECT1_0 = "NO";
    defparam add_20101_4.INJECT1_1 = "NO";
    CCU2D add_20101_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27205));
    defparam add_20101_2.INIT0 = 16'h1000;
    defparam add_20101_2.INIT1 = 16'h5555;
    defparam add_20101_2.INJECT1_0 = "NO";
    defparam add_20101_2.INJECT1_1 = "NO";
    FD1S3IX count_2643__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i0.GSR = "ENABLED";
    FD1S3AX clk_o_14 (.D(n8378), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2643__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i1.GSR = "ENABLED";
    FD1S3IX count_2643__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i2.GSR = "ENABLED";
    FD1S3IX count_2643__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i3.GSR = "ENABLED";
    FD1S3IX count_2643__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i4.GSR = "ENABLED";
    FD1S3IX count_2643__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i5.GSR = "ENABLED";
    FD1S3IX count_2643__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i6.GSR = "ENABLED";
    FD1S3IX count_2643__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i7.GSR = "ENABLED";
    FD1S3IX count_2643__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i8.GSR = "ENABLED";
    FD1S3IX count_2643__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i9.GSR = "ENABLED";
    FD1S3IX count_2643__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i10.GSR = "ENABLED";
    FD1S3IX count_2643__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i11.GSR = "ENABLED";
    FD1S3IX count_2643__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i12.GSR = "ENABLED";
    FD1S3IX count_2643__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i13.GSR = "ENABLED";
    FD1S3IX count_2643__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i14.GSR = "ENABLED";
    FD1S3IX count_2643__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i15.GSR = "ENABLED";
    FD1S3IX count_2643__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i16.GSR = "ENABLED";
    FD1S3IX count_2643__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i17.GSR = "ENABLED";
    FD1S3IX count_2643__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i18.GSR = "ENABLED";
    FD1S3IX count_2643__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i19.GSR = "ENABLED";
    FD1S3IX count_2643__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i20.GSR = "ENABLED";
    FD1S3IX count_2643__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i21.GSR = "ENABLED";
    FD1S3IX count_2643__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i22.GSR = "ENABLED";
    FD1S3IX count_2643__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i23.GSR = "ENABLED";
    FD1S3IX count_2643__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i24.GSR = "ENABLED";
    FD1S3IX count_2643__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i25.GSR = "ENABLED";
    FD1S3IX count_2643__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i26.GSR = "ENABLED";
    FD1S3IX count_2643__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i27.GSR = "ENABLED";
    FD1S3IX count_2643__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i28.GSR = "ENABLED";
    FD1S3IX count_2643__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i29.GSR = "ENABLED";
    FD1S3IX count_2643__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i30.GSR = "ENABLED";
    FD1S3IX count_2643__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16541), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2643__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000) 
//

module \ClockDividerP(factor=12000)  (GND_net, n8343, debug_c_c, n2954, 
            n30355, select_clk, n107) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n8343;
    input debug_c_c;
    input n2954;
    output n30355;
    output select_clk;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27256;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27255, n27254, n27253, n27252, n27251, n27250, n27249, 
        n27248, n27247, n27246, n27245, n27244, n27411;
    wire [31:0]n134;
    
    wire n27410, n27409, n27408, n27407, n27406, n27405, n27404, 
        n27403, n27402, n27401, n27400, n27399, n27398, n27397, 
        n27396, n28104, n15, n20, n16, n27, n40, n36, n28, 
        n18, n38, n32, n34, n24;
    
    CCU2D add_20100_28 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27256), 
          .S1(n8343));
    defparam add_20100_28.INIT0 = 16'h5555;
    defparam add_20100_28.INIT1 = 16'h0000;
    defparam add_20100_28.INJECT1_0 = "NO";
    defparam add_20100_28.INJECT1_1 = "NO";
    CCU2D add_20100_26 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27255), .COUT(n27256));
    defparam add_20100_26.INIT0 = 16'h5555;
    defparam add_20100_26.INIT1 = 16'h5555;
    defparam add_20100_26.INJECT1_0 = "NO";
    defparam add_20100_26.INJECT1_1 = "NO";
    CCU2D add_20100_24 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27254), .COUT(n27255));
    defparam add_20100_24.INIT0 = 16'h5555;
    defparam add_20100_24.INIT1 = 16'h5555;
    defparam add_20100_24.INJECT1_0 = "NO";
    defparam add_20100_24.INJECT1_1 = "NO";
    CCU2D add_20100_22 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27253), .COUT(n27254));
    defparam add_20100_22.INIT0 = 16'h5555;
    defparam add_20100_22.INIT1 = 16'h5555;
    defparam add_20100_22.INJECT1_0 = "NO";
    defparam add_20100_22.INJECT1_1 = "NO";
    CCU2D add_20100_20 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27252), .COUT(n27253));
    defparam add_20100_20.INIT0 = 16'h5555;
    defparam add_20100_20.INIT1 = 16'h5555;
    defparam add_20100_20.INJECT1_0 = "NO";
    defparam add_20100_20.INJECT1_1 = "NO";
    CCU2D add_20100_18 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27251), .COUT(n27252));
    defparam add_20100_18.INIT0 = 16'h5555;
    defparam add_20100_18.INIT1 = 16'h5555;
    defparam add_20100_18.INJECT1_0 = "NO";
    defparam add_20100_18.INJECT1_1 = "NO";
    CCU2D add_20100_16 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27250), .COUT(n27251));
    defparam add_20100_16.INIT0 = 16'h5555;
    defparam add_20100_16.INIT1 = 16'h5555;
    defparam add_20100_16.INJECT1_0 = "NO";
    defparam add_20100_16.INJECT1_1 = "NO";
    CCU2D add_20100_14 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27249), .COUT(n27250));
    defparam add_20100_14.INIT0 = 16'h5555;
    defparam add_20100_14.INIT1 = 16'h5555;
    defparam add_20100_14.INJECT1_0 = "NO";
    defparam add_20100_14.INJECT1_1 = "NO";
    CCU2D add_20100_12 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27248), .COUT(n27249));
    defparam add_20100_12.INIT0 = 16'h5555;
    defparam add_20100_12.INIT1 = 16'h5555;
    defparam add_20100_12.INJECT1_0 = "NO";
    defparam add_20100_12.INJECT1_1 = "NO";
    CCU2D add_20100_10 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27247), .COUT(n27248));
    defparam add_20100_10.INIT0 = 16'h5555;
    defparam add_20100_10.INIT1 = 16'h5555;
    defparam add_20100_10.INJECT1_0 = "NO";
    defparam add_20100_10.INJECT1_1 = "NO";
    CCU2D add_20100_8 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27246), .COUT(n27247));
    defparam add_20100_8.INIT0 = 16'h5555;
    defparam add_20100_8.INIT1 = 16'h5aaa;
    defparam add_20100_8.INJECT1_0 = "NO";
    defparam add_20100_8.INJECT1_1 = "NO";
    CCU2D add_20100_6 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27245), .COUT(n27246));
    defparam add_20100_6.INIT0 = 16'h5aaa;
    defparam add_20100_6.INIT1 = 16'h5aaa;
    defparam add_20100_6.INJECT1_0 = "NO";
    defparam add_20100_6.INJECT1_1 = "NO";
    CCU2D add_20100_4 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27244), 
          .COUT(n27245));
    defparam add_20100_4.INIT0 = 16'h5555;
    defparam add_20100_4.INIT1 = 16'h5aaa;
    defparam add_20100_4.INJECT1_0 = "NO";
    defparam add_20100_4.INJECT1_1 = "NO";
    CCU2D add_20100_2 (.A0(count[5]), .B0(count[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27244));
    defparam add_20100_2.INIT0 = 16'h7000;
    defparam add_20100_2.INIT1 = 16'h5aaa;
    defparam add_20100_2.INJECT1_0 = "NO";
    defparam add_20100_2.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27411), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_33.INIT1 = 16'h0000;
    defparam count_2642_add_4_33.INJECT1_0 = "NO";
    defparam count_2642_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27410), .COUT(n27411), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_31.INJECT1_0 = "NO";
    defparam count_2642_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27409), .COUT(n27410), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_29.INJECT1_0 = "NO";
    defparam count_2642_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27408), .COUT(n27409), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_27.INJECT1_0 = "NO";
    defparam count_2642_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27407), .COUT(n27408), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_25.INJECT1_0 = "NO";
    defparam count_2642_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27406), .COUT(n27407), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_23.INJECT1_0 = "NO";
    defparam count_2642_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27405), .COUT(n27406), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_21.INJECT1_0 = "NO";
    defparam count_2642_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27404), .COUT(n27405), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_19.INJECT1_0 = "NO";
    defparam count_2642_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27403), .COUT(n27404), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_17.INJECT1_0 = "NO";
    defparam count_2642_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27402), .COUT(n27403), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_15.INJECT1_0 = "NO";
    defparam count_2642_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27401), .COUT(n27402), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_13.INJECT1_0 = "NO";
    defparam count_2642_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27400), .COUT(n27401), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_11.INJECT1_0 = "NO";
    defparam count_2642_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27399), .COUT(n27400), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_9.INJECT1_0 = "NO";
    defparam count_2642_add_4_9.INJECT1_1 = "NO";
    FD1S3IX count_2642__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2954), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i0.GSR = "ENABLED";
    CCU2D count_2642_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27398), .COUT(n27399), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_7.INJECT1_0 = "NO";
    defparam count_2642_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27397), .COUT(n27398), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_5.INJECT1_0 = "NO";
    defparam count_2642_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27396), .COUT(n27397), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2642_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2642_add_4_3.INJECT1_0 = "NO";
    defparam count_2642_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2642_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27396), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642_add_4_1.INIT0 = 16'hF000;
    defparam count_2642_add_4_1.INIT1 = 16'h0555;
    defparam count_2642_add_4_1.INJECT1_0 = "NO";
    defparam count_2642_add_4_1.INJECT1_1 = "NO";
    LUT4 i23043_4_lut (.A(n28104), .B(n15), .C(n20), .D(n16), .Z(n30355)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i23043_4_lut.init = 16'h4000;
    LUT4 i20_4_lut (.A(n27), .B(n40), .C(n36), .D(n28), .Z(n28104)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[11]), .B(count[10]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(count[9]), .B(n18), .C(count[6]), .D(count[7]), 
         .Z(n20)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(count[1]), .B(count[4]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i6_2_lut (.A(count[28]), .B(count[12]), .Z(n27)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[5]), .B(n38), .C(n32), .D(count[20]), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(count[8]), .B(count[25]), .C(count[15]), .D(count[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[17]), .B(count[24]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i7_4_lut (.A(count[13]), .B(count[2]), .C(count[3]), .D(count[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i17_4_lut (.A(count[29]), .B(n34), .C(n24), .D(count[14]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(count[22]), .B(count[21]), .C(count[31]), .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(count[16]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[19]), .B(count[18]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    FD1S3AX clk_o_14 (.D(n107), .CK(debug_c_c), .Q(select_clk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=25, LSE_RCOL=48, LSE_LLINE=21, LSE_RLINE=23 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2642__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2954), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i1.GSR = "ENABLED";
    FD1S3IX count_2642__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2954), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i2.GSR = "ENABLED";
    FD1S3IX count_2642__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2954), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i3.GSR = "ENABLED";
    FD1S3IX count_2642__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2954), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i4.GSR = "ENABLED";
    FD1S3IX count_2642__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2954), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i5.GSR = "ENABLED";
    FD1S3IX count_2642__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2954), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i6.GSR = "ENABLED";
    FD1S3IX count_2642__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2954), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i7.GSR = "ENABLED";
    FD1S3IX count_2642__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2954), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i8.GSR = "ENABLED";
    FD1S3IX count_2642__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2954), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i9.GSR = "ENABLED";
    FD1S3IX count_2642__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i10.GSR = "ENABLED";
    FD1S3IX count_2642__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i11.GSR = "ENABLED";
    FD1S3IX count_2642__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i12.GSR = "ENABLED";
    FD1S3IX count_2642__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i13.GSR = "ENABLED";
    FD1S3IX count_2642__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i14.GSR = "ENABLED";
    FD1S3IX count_2642__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i15.GSR = "ENABLED";
    FD1S3IX count_2642__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i16.GSR = "ENABLED";
    FD1S3IX count_2642__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i17.GSR = "ENABLED";
    FD1S3IX count_2642__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i18.GSR = "ENABLED";
    FD1S3IX count_2642__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i19.GSR = "ENABLED";
    FD1S3IX count_2642__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i20.GSR = "ENABLED";
    FD1S3IX count_2642__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i21.GSR = "ENABLED";
    FD1S3IX count_2642__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i22.GSR = "ENABLED";
    FD1S3IX count_2642__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i23.GSR = "ENABLED";
    FD1S3IX count_2642__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i24.GSR = "ENABLED";
    FD1S3IX count_2642__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i25.GSR = "ENABLED";
    FD1S3IX count_2642__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i26.GSR = "ENABLED";
    FD1S3IX count_2642__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i27.GSR = "ENABLED";
    FD1S3IX count_2642__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i28.GSR = "ENABLED";
    FD1S3IX count_2642__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i29.GSR = "ENABLED";
    FD1S3IX count_2642__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i30.GSR = "ENABLED";
    FD1S3IX count_2642__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2954), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2642__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (debug_c_c, VCC_net, GND_net, 
            Stepper_Y_nFault_c, n31991, \read_size[0] , n13700, n96, 
            Stepper_Y_M0_c_0, n111, n579, prev_step_clk, step_clk, 
            limit_latched, prev_limit_latched, n14094, prev_select, 
            n31977, \register_addr[0] , \register_addr[1] , n27769, 
            n31953, databus, \div_factor_reg[9] , \div_factor_reg[6] , 
            \div_factor_reg[5] , \div_factor_reg[3] , \control_reg[7] , 
            n13667, n11927, Stepper_Y_En_c, Stepper_Y_Dir_c, \control_reg[3] , 
            Stepper_Y_M2_c_2, Stepper_Y_M1_c_1, \read_size[2] , n29768, 
            \steps_reg[9] , \steps_reg[6] , \steps_reg[5] , \steps_reg[3] , 
            n32, n29770, read_value, n4071, limit_c_1, n8476, n29788, 
            n31921, n21084, n21092, n6785, int_step, n22, n31919, 
            n31905, n16545, n7996, n8030) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    input n31991;
    output \read_size[0] ;
    input n13700;
    input n96;
    output Stepper_Y_M0_c_0;
    input n111;
    input n579;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    input n14094;
    output prev_select;
    input n31977;
    input \register_addr[0] ;
    input \register_addr[1] ;
    output n27769;
    input n31953;
    input [31:0]databus;
    output \div_factor_reg[9] ;
    output \div_factor_reg[6] ;
    output \div_factor_reg[5] ;
    output \div_factor_reg[3] ;
    output \control_reg[7] ;
    input n13667;
    input n11927;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output \control_reg[3] ;
    output Stepper_Y_M2_c_2;
    output Stepper_Y_M1_c_1;
    output \read_size[2] ;
    input n29768;
    output \steps_reg[9] ;
    output \steps_reg[6] ;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input n32;
    input n29770;
    output [31:0]read_value;
    input n4071;
    input limit_c_1;
    input n8476;
    input n29788;
    input n31921;
    input n21084;
    input n21092;
    input n6785;
    output int_step;
    input n22;
    input n31919;
    input n31905;
    input n16545;
    output n7996;
    output n8030;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire fault_latched;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n4072;
    
    wire n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n30338, n30339, n30340, n49, n62, n58, n50, n41, n60, 
        n54, n42, n27173;
    wire [31:0]n224;
    
    wire n27172;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n27171, n27170, n27169, n27168, n27167, n27166, n30311, 
        n30312, n30313, n27165, n27164, n27163, n27162, n27161, 
        n27160, n27159, n27158, n52, n38, n56, n46, n29780, 
        n29789, n29794, n29793, n29792, n29791, n29779, n29790, 
        n29771;
    wire [7:0]n8475;
    wire [31:0]n6720;
    
    wire n29777, n29787, n29786, n30266, n30267, n29785, n29784, 
        n29783;
    wire [31:0]n6756;
    
    wire n29782, n29778, n29776, n29775, n29774, n29772, n29773, 
        n29781, n30268;
    
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4072[0]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n96), .SP(n13700), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n111), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n14094), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31977), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i22928_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22928_3_lut.init = 16'hcaca;
    LUT4 i22929_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22929_3_lut.init = 16'hcaca;
    PFUMX i22930 (.BLUT(n30338), .ALUT(n30339), .C0(\register_addr[1] ), 
          .Z(n30340));
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27769)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27173), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27172), .COUT(n27173), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n31953), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n31953), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n31953), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n31953), .PD(n31991), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n31953), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n31953), .PD(n31991), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n31953), .PD(n31991), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n31953), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13667), .CD(n11927), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13667), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13667), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13667), .CD(n31991), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13667), .PD(n31991), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13667), .CD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13667), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27171), .COUT(n27172), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27170), .COUT(n27171), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27169), .COUT(n27170), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    FD1P3AX read_size__i2 (.D(n29768), .SP(n13700), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n4072[31]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4072[30]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4072[29]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4072[28]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4072[27]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4072[26]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4072[25]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4072[24]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4072[23]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4072[22]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4072[21]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4072[20]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4072[19]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4072[18]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4072[17]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4072[16]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4072[15]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4072[14]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4072[13]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4072[12]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4072[11]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4072[10]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4072[9]), .CK(debug_c_c), .CD(n31991), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4072[8]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4072[7]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4072[6]), .CK(debug_c_c), .CD(n31991), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4072[5]), .CK(debug_c_c), .CD(n31991), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4072[4]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4072[3]), .CK(debug_c_c), .CD(n31991), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4072[2]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4072[1]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27168), .COUT(n27169), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27167), .COUT(n27168), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27166), .COUT(n27167), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    PFUMX i22903 (.BLUT(n30311), .ALUT(n30312), .C0(\register_addr[0] ), 
          .Z(n30313));
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27165), .COUT(n27166), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27164), .COUT(n27165), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27163), .COUT(n27164), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27162), .COUT(n27163), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27161), .COUT(n27162), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27160), .COUT(n27161), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27159), .COUT(n27160), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27158), .COUT(n27159), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27158), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i1_4_lut (.A(div_factor_reg[31]), .B(n29770), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n29780)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_242 (.A(div_factor_reg[30]), .B(n29770), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29789)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_242.init = 16'hc088;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_243 (.A(div_factor_reg[29]), .B(n29770), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29794)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_243.init = 16'hc088;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_244 (.A(div_factor_reg[28]), .B(n29770), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n29793)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_244.init = 16'hc088;
    LUT4 i1_4_lut_adj_245 (.A(div_factor_reg[27]), .B(n29770), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n29792)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_245.init = 16'hc088;
    LUT4 i1_4_lut_adj_246 (.A(div_factor_reg[26]), .B(n29770), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n29791)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_246.init = 16'hc088;
    LUT4 i1_4_lut_adj_247 (.A(div_factor_reg[25]), .B(n29770), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n29779)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_247.init = 16'hc088;
    LUT4 i1_4_lut_adj_248 (.A(div_factor_reg[24]), .B(n29770), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n29790)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_248.init = 16'hc088;
    LUT4 i1_4_lut_adj_249 (.A(div_factor_reg[23]), .B(n29770), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n29771)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_249.init = 16'hc088;
    LUT4 i14792_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8475[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14792_2_lut.init = 16'h2222;
    LUT4 mux_1933_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n6720[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1933_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_250 (.A(div_factor_reg[22]), .B(n29770), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n29777)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_250.init = 16'hc088;
    LUT4 i1_4_lut_adj_251 (.A(div_factor_reg[21]), .B(n29770), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n29787)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_251.init = 16'hc088;
    LUT4 i1_4_lut_adj_252 (.A(div_factor_reg[20]), .B(n29770), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n29786)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_252.init = 16'hc088;
    LUT4 i22856_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22856_3_lut.init = 16'hcaca;
    LUT4 i22857_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22857_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i31 (.D(n29780), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29789), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29794), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29793), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29792), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29791), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29779), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29790), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29771), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    LUT4 mux_1933_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6720[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1933_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_253 (.A(div_factor_reg[19]), .B(n29770), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n29785)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_253.init = 16'hc088;
    LUT4 i1_4_lut_adj_254 (.A(div_factor_reg[18]), .B(n29770), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n29784)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_254.init = 16'hc088;
    LUT4 i1_4_lut_adj_255 (.A(div_factor_reg[17]), .B(n29770), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n29783)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_255.init = 16'hc088;
    PFUMX mux_1937_i5 (.BLUT(n8475[4]), .ALUT(n6720[4]), .C0(\register_addr[1] ), 
          .Z(n6756[4]));
    LUT4 mux_1582_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4071), .Z(n4072[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_256 (.A(div_factor_reg[16]), .B(n29770), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n29782)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_256.init = 16'hc088;
    LUT4 i1_4_lut_adj_257 (.A(div_factor_reg[15]), .B(n29770), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n29778)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_257.init = 16'hc088;
    LUT4 i1_4_lut_adj_258 (.A(div_factor_reg[14]), .B(n29770), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n29776)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_258.init = 16'hc088;
    LUT4 i1_4_lut_adj_259 (.A(div_factor_reg[13]), .B(n29770), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n29775)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_259.init = 16'hc088;
    FD1P3AX read_value__i22 (.D(n29777), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29787), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_260 (.A(div_factor_reg[12]), .B(n29770), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n29774)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_260.init = 16'hc088;
    LUT4 i1_4_lut_adj_261 (.A(div_factor_reg[11]), .B(n29770), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n29772)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_261.init = 16'hc088;
    LUT4 i1_4_lut_adj_262 (.A(div_factor_reg[10]), .B(n29770), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n29773)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_262.init = 16'hc088;
    LUT4 i1_4_lut_adj_263 (.A(div_factor_reg[8]), .B(n29770), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29781)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_263.init = 16'hc088;
    FD1P3AX read_value__i20 (.D(n29786), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    PFUMX i22858 (.BLUT(n30266), .ALUT(n30267), .C0(\register_addr[1] ), 
          .Z(n30268));
    LUT4 mux_1582_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4071), 
         .Z(n4072[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4071), 
         .Z(n4072[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i31_3_lut.init = 16'hcaca;
    PFUMX mux_1937_i8 (.BLUT(n8476), .ALUT(n6720[7]), .C0(\register_addr[1] ), 
          .Z(n6756[7]));
    LUT4 mux_1582_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4071), 
         .Z(n4072[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4071), 
         .Z(n4072[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4071), 
         .Z(n4072[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i28_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i19 (.D(n29785), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29784), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29783), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29782), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29778), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29776), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29775), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29774), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29772), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29773), .SP(n13700), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29788), .SP(n13700), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29781), .SP(n13700), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6756[7]), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n21084), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n21092), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6756[4]), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6785), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30313), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30268), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1582_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4071), 
         .Z(n4072[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4071), 
         .Z(n4072[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4071), 
         .Z(n4072[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4071), 
         .Z(n4072[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i24_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n31919), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1582_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4071), 
         .Z(n4072[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i23_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n30340), .SP(n13700), .CD(n31921), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=599, LSE_RLINE=612 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_1582_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4071), 
         .Z(n4072[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4071), 
         .Z(n4072[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4071), 
         .Z(n4072[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4071), 
         .Z(n4072[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4071), 
         .Z(n4072[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4071), 
         .Z(n4072[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4071), 
         .Z(n4072[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4071), 
         .Z(n4072[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4071), 
         .Z(n4072[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4071), 
         .Z(n4072[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4071), 
         .Z(n4072[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4071), 
         .Z(n4072[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4071), .Z(n4072[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4071), .Z(n4072[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4071), .Z(n4072[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4071), .Z(n4072[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4071), .Z(n4072[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4071), .Z(n4072[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4071), .Z(n4072[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4071), .Z(n4072[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4071), .Z(n4072[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1582_i2_3_lut.init = 16'hcaca;
    LUT4 i22901_3_lut (.A(Stepper_Y_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22901_3_lut.init = 16'hcaca;
    LUT4 i22902_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22902_3_lut.init = 16'hcaca;
    ClockDivider_U7 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n31991(n31991), .n31905(n31905), .n16545(n16545), 
            .div_factor_reg({div_factor_reg[31:10], \div_factor_reg[9] , 
            div_factor_reg[8:7], \div_factor_reg[6] , \div_factor_reg[5] , 
            div_factor_reg[4], \div_factor_reg[3] , div_factor_reg[2:0]}), 
            .n7996(n7996), .n8030(n8030)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (GND_net, step_clk, debug_c_c, n31991, n31905, 
            n16545, div_factor_reg, n7996, n8030) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31991;
    input n31905;
    input n16545;
    input [31:0]div_factor_reg;
    output n7996;
    output n8030;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27243;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27242, n27241, n27240, n27239, n27238, n27237, n27236, 
        n27235, n27234, n27233, n27232, n27231, n27230, n27229, 
        n27228, n7961, n26957, n26956;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26955, n26954, n26953, n26952, n26951, n26950, n26949, 
        n26948, n26947, n26946, n26945, n26944, n26943, n26942, 
        n26941;
    wire [31:0]n40;
    
    wire n26940, n26939, n26938, n26937, n26936, n26935, n26934, 
        n26933, n26932, n26931, n26930, n26929, n26928, n26927, 
        n26926, n26925, n26924, n26923, n26922, n26921, n26920, 
        n27109, n26919, n26918, n27108, n27107, n27106, n27105, 
        n26917, n27104, n27103, n27102, n27101, n26916, n26915, 
        n26914, n26913, n27100, n27099, n26912, n26911, n27098, 
        n27097, n27096, n26910, n27095, n27094;
    
    CCU2D count_2637_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27243), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_33.INIT1 = 16'h0000;
    defparam count_2637_add_4_33.INJECT1_0 = "NO";
    defparam count_2637_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27242), .COUT(n27243), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_31.INJECT1_0 = "NO";
    defparam count_2637_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27241), .COUT(n27242), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_29.INJECT1_0 = "NO";
    defparam count_2637_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27240), .COUT(n27241), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_27.INJECT1_0 = "NO";
    defparam count_2637_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27239), .COUT(n27240), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_25.INJECT1_0 = "NO";
    defparam count_2637_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27238), .COUT(n27239), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_23.INJECT1_0 = "NO";
    defparam count_2637_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27237), .COUT(n27238), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_21.INJECT1_0 = "NO";
    defparam count_2637_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27236), .COUT(n27237), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_19.INJECT1_0 = "NO";
    defparam count_2637_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27235), .COUT(n27236), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_17.INJECT1_0 = "NO";
    defparam count_2637_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27234), .COUT(n27235), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_15.INJECT1_0 = "NO";
    defparam count_2637_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27233), .COUT(n27234), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_13.INJECT1_0 = "NO";
    defparam count_2637_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27232), .COUT(n27233), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_11.INJECT1_0 = "NO";
    defparam count_2637_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27231), .COUT(n27232), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_9.INJECT1_0 = "NO";
    defparam count_2637_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27230), .COUT(n27231), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_7.INJECT1_0 = "NO";
    defparam count_2637_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27229), .COUT(n27230), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_5.INJECT1_0 = "NO";
    defparam count_2637_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27228), .COUT(n27229), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2637_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2637_add_4_3.INJECT1_0 = "NO";
    defparam count_2637_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2637_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27228), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637_add_4_1.INIT0 = 16'hF000;
    defparam count_2637_add_4_1.INIT1 = 16'h0555;
    defparam count_2637_add_4_1.INJECT1_0 = "NO";
    defparam count_2637_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7961), .CK(debug_c_c), .CD(n31991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2039_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26957), .S1(n7961));
    defparam sub_2039_add_2_33.INIT0 = 16'h5555;
    defparam sub_2039_add_2_33.INIT1 = 16'h0000;
    defparam sub_2039_add_2_33.INJECT1_0 = "NO";
    defparam sub_2039_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26956), .COUT(n26957));
    defparam sub_2039_add_2_31.INIT0 = 16'h5999;
    defparam sub_2039_add_2_31.INIT1 = 16'h5999;
    defparam sub_2039_add_2_31.INJECT1_0 = "NO";
    defparam sub_2039_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26955), .COUT(n26956));
    defparam sub_2039_add_2_29.INIT0 = 16'h5999;
    defparam sub_2039_add_2_29.INIT1 = 16'h5999;
    defparam sub_2039_add_2_29.INJECT1_0 = "NO";
    defparam sub_2039_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26954), .COUT(n26955));
    defparam sub_2039_add_2_27.INIT0 = 16'h5999;
    defparam sub_2039_add_2_27.INIT1 = 16'h5999;
    defparam sub_2039_add_2_27.INJECT1_0 = "NO";
    defparam sub_2039_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26953), .COUT(n26954));
    defparam sub_2039_add_2_25.INIT0 = 16'h5999;
    defparam sub_2039_add_2_25.INIT1 = 16'h5999;
    defparam sub_2039_add_2_25.INJECT1_0 = "NO";
    defparam sub_2039_add_2_25.INJECT1_1 = "NO";
    FD1S3IX count_2637__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i0.GSR = "ENABLED";
    CCU2D sub_2039_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26952), .COUT(n26953));
    defparam sub_2039_add_2_23.INIT0 = 16'h5999;
    defparam sub_2039_add_2_23.INIT1 = 16'h5999;
    defparam sub_2039_add_2_23.INJECT1_0 = "NO";
    defparam sub_2039_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26951), .COUT(n26952));
    defparam sub_2039_add_2_21.INIT0 = 16'h5999;
    defparam sub_2039_add_2_21.INIT1 = 16'h5999;
    defparam sub_2039_add_2_21.INJECT1_0 = "NO";
    defparam sub_2039_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26950), .COUT(n26951));
    defparam sub_2039_add_2_19.INIT0 = 16'h5999;
    defparam sub_2039_add_2_19.INIT1 = 16'h5999;
    defparam sub_2039_add_2_19.INJECT1_0 = "NO";
    defparam sub_2039_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26949), .COUT(n26950));
    defparam sub_2039_add_2_17.INIT0 = 16'h5999;
    defparam sub_2039_add_2_17.INIT1 = 16'h5999;
    defparam sub_2039_add_2_17.INJECT1_0 = "NO";
    defparam sub_2039_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26948), .COUT(n26949));
    defparam sub_2039_add_2_15.INIT0 = 16'h5999;
    defparam sub_2039_add_2_15.INIT1 = 16'h5999;
    defparam sub_2039_add_2_15.INJECT1_0 = "NO";
    defparam sub_2039_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26947), .COUT(n26948));
    defparam sub_2039_add_2_13.INIT0 = 16'h5999;
    defparam sub_2039_add_2_13.INIT1 = 16'h5999;
    defparam sub_2039_add_2_13.INJECT1_0 = "NO";
    defparam sub_2039_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26946), .COUT(n26947));
    defparam sub_2039_add_2_11.INIT0 = 16'h5999;
    defparam sub_2039_add_2_11.INIT1 = 16'h5999;
    defparam sub_2039_add_2_11.INJECT1_0 = "NO";
    defparam sub_2039_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26945), .COUT(n26946));
    defparam sub_2039_add_2_9.INIT0 = 16'h5999;
    defparam sub_2039_add_2_9.INIT1 = 16'h5999;
    defparam sub_2039_add_2_9.INJECT1_0 = "NO";
    defparam sub_2039_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26944), .COUT(n26945));
    defparam sub_2039_add_2_7.INIT0 = 16'h5999;
    defparam sub_2039_add_2_7.INIT1 = 16'h5999;
    defparam sub_2039_add_2_7.INJECT1_0 = "NO";
    defparam sub_2039_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26943), .COUT(n26944));
    defparam sub_2039_add_2_5.INIT0 = 16'h5999;
    defparam sub_2039_add_2_5.INIT1 = 16'h5999;
    defparam sub_2039_add_2_5.INJECT1_0 = "NO";
    defparam sub_2039_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26942), .COUT(n26943));
    defparam sub_2039_add_2_3.INIT0 = 16'h5999;
    defparam sub_2039_add_2_3.INIT1 = 16'h5999;
    defparam sub_2039_add_2_3.INJECT1_0 = "NO";
    defparam sub_2039_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2039_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26942));
    defparam sub_2039_add_2_1.INIT0 = 16'h0000;
    defparam sub_2039_add_2_1.INIT1 = 16'h5999;
    defparam sub_2039_add_2_1.INJECT1_0 = "NO";
    defparam sub_2039_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2041_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26941), .S1(n7996));
    defparam sub_2041_add_2_33.INIT0 = 16'h5999;
    defparam sub_2041_add_2_33.INIT1 = 16'h0000;
    defparam sub_2041_add_2_33.INJECT1_0 = "NO";
    defparam sub_2041_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26940), .COUT(n26941));
    defparam sub_2041_add_2_31.INIT0 = 16'h5999;
    defparam sub_2041_add_2_31.INIT1 = 16'h5999;
    defparam sub_2041_add_2_31.INJECT1_0 = "NO";
    defparam sub_2041_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26939), .COUT(n26940));
    defparam sub_2041_add_2_29.INIT0 = 16'h5999;
    defparam sub_2041_add_2_29.INIT1 = 16'h5999;
    defparam sub_2041_add_2_29.INJECT1_0 = "NO";
    defparam sub_2041_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26938), .COUT(n26939));
    defparam sub_2041_add_2_27.INIT0 = 16'h5999;
    defparam sub_2041_add_2_27.INIT1 = 16'h5999;
    defparam sub_2041_add_2_27.INJECT1_0 = "NO";
    defparam sub_2041_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26937), .COUT(n26938));
    defparam sub_2041_add_2_25.INIT0 = 16'h5999;
    defparam sub_2041_add_2_25.INIT1 = 16'h5999;
    defparam sub_2041_add_2_25.INJECT1_0 = "NO";
    defparam sub_2041_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26936), .COUT(n26937));
    defparam sub_2041_add_2_23.INIT0 = 16'h5999;
    defparam sub_2041_add_2_23.INIT1 = 16'h5999;
    defparam sub_2041_add_2_23.INJECT1_0 = "NO";
    defparam sub_2041_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26935), .COUT(n26936));
    defparam sub_2041_add_2_21.INIT0 = 16'h5999;
    defparam sub_2041_add_2_21.INIT1 = 16'h5999;
    defparam sub_2041_add_2_21.INJECT1_0 = "NO";
    defparam sub_2041_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26934), .COUT(n26935));
    defparam sub_2041_add_2_19.INIT0 = 16'h5999;
    defparam sub_2041_add_2_19.INIT1 = 16'h5999;
    defparam sub_2041_add_2_19.INJECT1_0 = "NO";
    defparam sub_2041_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26933), .COUT(n26934));
    defparam sub_2041_add_2_17.INIT0 = 16'h5999;
    defparam sub_2041_add_2_17.INIT1 = 16'h5999;
    defparam sub_2041_add_2_17.INJECT1_0 = "NO";
    defparam sub_2041_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26932), .COUT(n26933));
    defparam sub_2041_add_2_15.INIT0 = 16'h5999;
    defparam sub_2041_add_2_15.INIT1 = 16'h5999;
    defparam sub_2041_add_2_15.INJECT1_0 = "NO";
    defparam sub_2041_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26931), .COUT(n26932));
    defparam sub_2041_add_2_13.INIT0 = 16'h5999;
    defparam sub_2041_add_2_13.INIT1 = 16'h5999;
    defparam sub_2041_add_2_13.INJECT1_0 = "NO";
    defparam sub_2041_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26930), .COUT(n26931));
    defparam sub_2041_add_2_11.INIT0 = 16'h5999;
    defparam sub_2041_add_2_11.INIT1 = 16'h5999;
    defparam sub_2041_add_2_11.INJECT1_0 = "NO";
    defparam sub_2041_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26929), .COUT(n26930));
    defparam sub_2041_add_2_9.INIT0 = 16'h5999;
    defparam sub_2041_add_2_9.INIT1 = 16'h5999;
    defparam sub_2041_add_2_9.INJECT1_0 = "NO";
    defparam sub_2041_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26928), .COUT(n26929));
    defparam sub_2041_add_2_7.INIT0 = 16'h5999;
    defparam sub_2041_add_2_7.INIT1 = 16'h5999;
    defparam sub_2041_add_2_7.INJECT1_0 = "NO";
    defparam sub_2041_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26927), .COUT(n26928));
    defparam sub_2041_add_2_5.INIT0 = 16'h5999;
    defparam sub_2041_add_2_5.INIT1 = 16'h5999;
    defparam sub_2041_add_2_5.INJECT1_0 = "NO";
    defparam sub_2041_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2041_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26926), .COUT(n26927));
    defparam sub_2041_add_2_3.INIT0 = 16'h5999;
    defparam sub_2041_add_2_3.INIT1 = 16'h5999;
    defparam sub_2041_add_2_3.INJECT1_0 = "NO";
    defparam sub_2041_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31905), .CD(n16545), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31905), .PD(n16545), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2041_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26926));
    defparam sub_2041_add_2_1.INIT0 = 16'h0000;
    defparam sub_2041_add_2_1.INIT1 = 16'h5999;
    defparam sub_2041_add_2_1.INJECT1_0 = "NO";
    defparam sub_2041_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26925), .S1(n8030));
    defparam sub_2042_add_2_33.INIT0 = 16'hf555;
    defparam sub_2042_add_2_33.INIT1 = 16'h0000;
    defparam sub_2042_add_2_33.INJECT1_0 = "NO";
    defparam sub_2042_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26924), .COUT(n26925));
    defparam sub_2042_add_2_31.INIT0 = 16'hf555;
    defparam sub_2042_add_2_31.INIT1 = 16'hf555;
    defparam sub_2042_add_2_31.INJECT1_0 = "NO";
    defparam sub_2042_add_2_31.INJECT1_1 = "NO";
    FD1S3IX count_2637__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i1.GSR = "ENABLED";
    FD1S3IX count_2637__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i2.GSR = "ENABLED";
    FD1S3IX count_2637__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i3.GSR = "ENABLED";
    FD1S3IX count_2637__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i4.GSR = "ENABLED";
    FD1S3IX count_2637__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i5.GSR = "ENABLED";
    FD1S3IX count_2637__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i6.GSR = "ENABLED";
    FD1S3IX count_2637__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i7.GSR = "ENABLED";
    FD1S3IX count_2637__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i8.GSR = "ENABLED";
    FD1S3IX count_2637__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i9.GSR = "ENABLED";
    FD1S3IX count_2637__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i10.GSR = "ENABLED";
    FD1S3IX count_2637__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i11.GSR = "ENABLED";
    FD1S3IX count_2637__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i12.GSR = "ENABLED";
    FD1S3IX count_2637__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i13.GSR = "ENABLED";
    FD1S3IX count_2637__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i14.GSR = "ENABLED";
    FD1S3IX count_2637__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i15.GSR = "ENABLED";
    FD1S3IX count_2637__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i16.GSR = "ENABLED";
    FD1S3IX count_2637__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i17.GSR = "ENABLED";
    FD1S3IX count_2637__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i18.GSR = "ENABLED";
    FD1S3IX count_2637__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i19.GSR = "ENABLED";
    FD1S3IX count_2637__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i20.GSR = "ENABLED";
    FD1S3IX count_2637__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i21.GSR = "ENABLED";
    FD1S3IX count_2637__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i22.GSR = "ENABLED";
    FD1S3IX count_2637__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i23.GSR = "ENABLED";
    FD1S3IX count_2637__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i24.GSR = "ENABLED";
    FD1S3IX count_2637__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i25.GSR = "ENABLED";
    FD1S3IX count_2637__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i26.GSR = "ENABLED";
    FD1S3IX count_2637__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i27.GSR = "ENABLED";
    FD1S3IX count_2637__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i28.GSR = "ENABLED";
    FD1S3IX count_2637__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i29.GSR = "ENABLED";
    FD1S3IX count_2637__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i30.GSR = "ENABLED";
    FD1S3IX count_2637__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31905), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2637__i31.GSR = "ENABLED";
    CCU2D sub_2042_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26923), .COUT(n26924));
    defparam sub_2042_add_2_29.INIT0 = 16'hf555;
    defparam sub_2042_add_2_29.INIT1 = 16'hf555;
    defparam sub_2042_add_2_29.INJECT1_0 = "NO";
    defparam sub_2042_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26922), .COUT(n26923));
    defparam sub_2042_add_2_27.INIT0 = 16'hf555;
    defparam sub_2042_add_2_27.INIT1 = 16'hf555;
    defparam sub_2042_add_2_27.INJECT1_0 = "NO";
    defparam sub_2042_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26921), .COUT(n26922));
    defparam sub_2042_add_2_25.INIT0 = 16'hf555;
    defparam sub_2042_add_2_25.INIT1 = 16'hf555;
    defparam sub_2042_add_2_25.INJECT1_0 = "NO";
    defparam sub_2042_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26920), .COUT(n26921));
    defparam sub_2042_add_2_23.INIT0 = 16'hf555;
    defparam sub_2042_add_2_23.INIT1 = 16'hf555;
    defparam sub_2042_add_2_23.INJECT1_0 = "NO";
    defparam sub_2042_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27109), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26919), .COUT(n26920));
    defparam sub_2042_add_2_21.INIT0 = 16'hf555;
    defparam sub_2042_add_2_21.INIT1 = 16'hf555;
    defparam sub_2042_add_2_21.INJECT1_0 = "NO";
    defparam sub_2042_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26918), .COUT(n26919));
    defparam sub_2042_add_2_19.INIT0 = 16'hf555;
    defparam sub_2042_add_2_19.INIT1 = 16'hf555;
    defparam sub_2042_add_2_19.INJECT1_0 = "NO";
    defparam sub_2042_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27108), .COUT(n27109), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27107), .COUT(n27108), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27106), .COUT(n27107), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27105), .COUT(n27106), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26917), .COUT(n26918));
    defparam sub_2042_add_2_17.INIT0 = 16'hf555;
    defparam sub_2042_add_2_17.INIT1 = 16'hf555;
    defparam sub_2042_add_2_17.INJECT1_0 = "NO";
    defparam sub_2042_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27104), .COUT(n27105), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27103), .COUT(n27104), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27102), .COUT(n27103), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27101), .COUT(n27102), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26916), .COUT(n26917));
    defparam sub_2042_add_2_15.INIT0 = 16'hf555;
    defparam sub_2042_add_2_15.INIT1 = 16'hf555;
    defparam sub_2042_add_2_15.INJECT1_0 = "NO";
    defparam sub_2042_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26915), .COUT(n26916));
    defparam sub_2042_add_2_13.INIT0 = 16'hf555;
    defparam sub_2042_add_2_13.INIT1 = 16'hf555;
    defparam sub_2042_add_2_13.INJECT1_0 = "NO";
    defparam sub_2042_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26914), .COUT(n26915));
    defparam sub_2042_add_2_11.INIT0 = 16'hf555;
    defparam sub_2042_add_2_11.INIT1 = 16'hf555;
    defparam sub_2042_add_2_11.INJECT1_0 = "NO";
    defparam sub_2042_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26913), .COUT(n26914));
    defparam sub_2042_add_2_9.INIT0 = 16'hf555;
    defparam sub_2042_add_2_9.INIT1 = 16'hf555;
    defparam sub_2042_add_2_9.INJECT1_0 = "NO";
    defparam sub_2042_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27100), .COUT(n27101), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27099), .COUT(n27100), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26912), .COUT(n26913));
    defparam sub_2042_add_2_7.INIT0 = 16'hf555;
    defparam sub_2042_add_2_7.INIT1 = 16'hf555;
    defparam sub_2042_add_2_7.INJECT1_0 = "NO";
    defparam sub_2042_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26911), .COUT(n26912));
    defparam sub_2042_add_2_5.INIT0 = 16'hf555;
    defparam sub_2042_add_2_5.INIT1 = 16'hf555;
    defparam sub_2042_add_2_5.INJECT1_0 = "NO";
    defparam sub_2042_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27098), .COUT(n27099), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27097), .COUT(n27098), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27096), .COUT(n27097), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26910), .COUT(n26911));
    defparam sub_2042_add_2_3.INIT0 = 16'hf555;
    defparam sub_2042_add_2_3.INIT1 = 16'hf555;
    defparam sub_2042_add_2_3.INJECT1_0 = "NO";
    defparam sub_2042_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27095), .COUT(n27096), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27094), .COUT(n27095), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27094), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2042_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26910));
    defparam sub_2042_add_2_1.INIT0 = 16'h0000;
    defparam sub_2042_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2042_add_2_1.INJECT1_0 = "NO";
    defparam sub_2042_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (read_value, debug_c_c, n2850, 
            n31991, n3899, VCC_net, GND_net, Stepper_A_nFault_c, \read_size[0] , 
            n29798, Stepper_A_M0_c_0, n22330, n579, limit_latched, 
            prev_limit_latched, n14661, prev_select, n31938, n32, 
            n32_adj_37, prev_step_clk, step_clk, n31918, n22, n32_adj_38, 
            prev_step_clk_adj_39, step_clk_adj_40, n31919, n22_adj_41, 
            prev_step_clk_adj_42, n34, step_clk_adj_43, n31920, n24, 
            \register_addr[1] , \register_addr[0] , \read_size[2] , n94, 
            Stepper_A_M1_c_1, n13710, \databus[1] , Stepper_A_M2_c_2, 
            \databus[2] , \databus[3] , \databus[4] , Stepper_A_Dir_c, 
            \databus[5] , Stepper_A_En_c, \databus[6] , \control_reg[7] , 
            n11981, \databus[7] , n31910, \databus[8] , \databus[9] , 
            \databus[10] , \databus[11] , \databus[12] , \databus[13] , 
            \databus[14] , \databus[15] , \databus[16] , \databus[17] , 
            \databus[18] , \databus[19] , \databus[20] , \databus[21] , 
            \databus[22] , \databus[23] , \databus[24] , \databus[25] , 
            \databus[26] , \databus[27] , \databus[28] , \databus[29] , 
            \databus[30] , \databus[31] , n224, n31911, n32056, n13323, 
            n32003, n30489, limit_c_3, n27766, Stepper_A_Step_c, n8494, 
            n31903, n16566, n8204, n8238) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2850;
    input n31991;
    input [31:0]n3899;
    input VCC_net;
    input GND_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n29798;
    output Stepper_A_M0_c_0;
    input n22330;
    input n579;
    output limit_latched;
    output prev_limit_latched;
    input n14661;
    output prev_select;
    input n31938;
    input n32;
    input n32_adj_37;
    input prev_step_clk;
    input step_clk;
    output n31918;
    output n22;
    input n32_adj_38;
    input prev_step_clk_adj_39;
    input step_clk_adj_40;
    output n31919;
    output n22_adj_41;
    input prev_step_clk_adj_42;
    input n34;
    input step_clk_adj_43;
    output n31920;
    output n24;
    input \register_addr[1] ;
    input \register_addr[0] ;
    output \read_size[2] ;
    input n94;
    output Stepper_A_M1_c_1;
    input n13710;
    input \databus[1] ;
    output Stepper_A_M2_c_2;
    input \databus[2] ;
    input \databus[3] ;
    input \databus[4] ;
    output Stepper_A_Dir_c;
    input \databus[5] ;
    output Stepper_A_En_c;
    input \databus[6] ;
    output \control_reg[7] ;
    input n11981;
    input \databus[7] ;
    input n31910;
    input \databus[8] ;
    input \databus[9] ;
    input \databus[10] ;
    input \databus[11] ;
    input \databus[12] ;
    input \databus[13] ;
    input \databus[14] ;
    input \databus[15] ;
    input \databus[16] ;
    input \databus[17] ;
    input \databus[18] ;
    input \databus[19] ;
    input \databus[20] ;
    input \databus[21] ;
    input \databus[22] ;
    input \databus[23] ;
    input \databus[24] ;
    input \databus[25] ;
    input \databus[26] ;
    input \databus[27] ;
    input \databus[28] ;
    input \databus[29] ;
    input \databus[30] ;
    input \databus[31] ;
    output [31:0]n224;
    input n31911;
    input n32056;
    input n13323;
    input n32003;
    output n30489;
    input limit_c_3;
    output n27766;
    output Stepper_A_Step_c;
    input n8494;
    input n31903;
    input n16566;
    output n8204;
    output n8238;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n30262;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire fault_latched, prev_step_clk_c, step_clk_c, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n31917, n22_c;
    wire [31:0]n100;
    
    wire n30310, n30265, n30308, n30309;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [7:0]n8493;
    wire [31:0]n7348;
    
    wire n27141, n27140, n27139, n27138, n27137, n27136, n27135, 
        n27134, n27133, n27132, n27131, n27130, n27129, n27128, 
        n27127, n27126, n30260, n30261, n30263, n30264, int_step, 
        n49, n62_adj_131, n58_adj_132, n50_adj_133, n41, n60_adj_134, 
        n54_adj_135, n42_adj_136, n52_adj_137, n38_adj_138, n56_adj_139, 
        n46_adj_140;
    
    FD1P3AX read_value__i0 (.D(n30262), .SP(n2850), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3899[0]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n29798), .SP(n2850), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n22330), .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk_c), .CK(debug_c_c), .Q(prev_step_clk_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n14661), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31938), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_300 (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .Z(n31917)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_300.init = 16'h2020;
    LUT4 i1_4_lut_4_lut (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .D(n31991), .Z(n22_c)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut.init = 16'h002c;
    LUT4 i2_3_lut_rep_301 (.A(n32_adj_37), .B(prev_step_clk), .C(step_clk), 
         .Z(n31918)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_301.init = 16'h2020;
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_239 (.A(n32_adj_37), .B(prev_step_clk), .C(step_clk), 
         .D(n31991), .Z(n22)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_239.init = 16'h002c;
    LUT4 i2_3_lut_rep_302 (.A(n32_adj_38), .B(prev_step_clk_adj_39), .C(step_clk_adj_40), 
         .Z(n31919)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_302.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_adj_240 (.A(n32_adj_38), .B(prev_step_clk_adj_39), 
         .C(step_clk_adj_40), .D(n31991), .Z(n22_adj_41)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_240.init = 16'h002c;
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30310), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30265), .SP(n2850), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_303 (.A(prev_step_clk_adj_42), .B(n34), .C(step_clk_adj_43), 
         .Z(n31920)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_303.init = 16'h4040;
    LUT4 i1_4_lut_4_lut_adj_241 (.A(prev_step_clk_adj_42), .B(n34), .C(step_clk_adj_43), 
         .D(n31991), .Z(n24)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_241.init = 16'h004a;
    LUT4 i14760_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14760_4_lut.init = 16'hc088;
    LUT4 i14761_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14761_4_lut.init = 16'hc088;
    PFUMX i22900 (.BLUT(n30308), .ALUT(n30309), .C0(\register_addr[0] ), 
          .Z(n30310));
    FD1S3IX steps_reg__i1 (.D(n3899[1]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3899[2]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3899[3]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3899[4]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3899[5]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3899[6]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3899[7]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3899[8]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3899[9]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3899[10]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3899[11]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3899[12]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3899[13]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3899[14]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3899[15]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3899[16]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3899[17]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3899[18]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3899[19]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3899[20]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3899[21]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3899[22]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3899[23]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3899[24]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3899[25]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3899[26]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3899[27]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3899[28]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3899[29]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3899[30]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3899[31]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n94), .SP(n2850), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(\databus[1] ), .SP(n13710), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(\databus[2] ), .SP(n13710), .CD(n31991), 
            .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(\databus[3] ), .SP(n13710), .PD(n31991), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(\databus[4] ), .SP(n13710), .CD(n31991), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(\databus[5] ), .SP(n13710), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(\databus[6] ), .SP(n13710), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(\databus[7] ), .SP(n13710), .CD(n11981), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(\databus[1] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(\databus[2] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(\databus[3] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(\databus[4] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(\databus[5] ), .SP(n31910), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(\databus[6] ), .SP(n31910), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(\databus[7] ), .SP(n31910), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(\databus[8] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(\databus[9] ), .SP(n31910), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(\databus[10] ), .SP(n31910), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(\databus[11] ), .SP(n31910), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(\databus[12] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(\databus[13] ), .SP(n31910), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(\databus[14] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(\databus[15] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(\databus[16] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(\databus[17] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(\databus[18] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(\databus[19] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(\databus[20] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(\databus[21] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(\databus[22] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(\databus[23] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(\databus[24] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(\databus[25] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(\databus[26] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(\databus[27] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(\databus[28] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(\databus[29] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(\databus[30] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(\databus[31] ), .SP(n31910), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=629, LSE_RLINE=642 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i14762_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14762_4_lut.init = 16'hc088;
    LUT4 i14749_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8493[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14749_2_lut.init = 16'h2222;
    LUT4 mux_1985_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7348[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1985_i4_3_lut.init = 16'hcaca;
    LUT4 i14763_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14763_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27141), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27140), .COUT(n27141), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    LUT4 i14748_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8493[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14748_2_lut.init = 16'h2222;
    LUT4 mux_1985_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7348[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1985_i5_3_lut.init = 16'hcaca;
    LUT4 i14747_2_lut (.A(Stepper_A_Dir_c), .B(\register_addr[0] ), .Z(n8493[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14747_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27139), .COUT(n27140), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27138), .COUT(n27139), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    LUT4 mux_1985_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7348[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1985_i6_3_lut.init = 16'hcaca;
    LUT4 i14764_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14764_4_lut.init = 16'hc088;
    LUT4 i14746_2_lut (.A(Stepper_A_En_c), .B(\register_addr[0] ), .Z(n8493[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14746_2_lut.init = 16'h2222;
    LUT4 i14765_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14765_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27137), .COUT(n27138), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    LUT4 i14766_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14766_4_lut.init = 16'hc088;
    LUT4 mux_1985_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7348[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1985_i7_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27136), .COUT(n27137), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    LUT4 mux_1985_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n7348[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1985_i8_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27135), .COUT(n27136), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27134), .COUT(n27135), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27133), .COUT(n27134), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27132), .COUT(n27133), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27131), .COUT(n27132), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27130), .COUT(n27131), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27129), .COUT(n27130), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27128), .COUT(n27129), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27127), .COUT(n27128), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 i14767_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14767_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27126), .COUT(n27127), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk_c), .D1(prev_step_clk_c), 
          .COUT(n27126), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i22850_3_lut (.A(Stepper_A_M0_c_0), .B(div_factor_reg[0]), .C(\register_addr[1] ), 
         .Z(n30260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22850_3_lut.init = 16'hcaca;
    LUT4 i22851_3_lut (.A(limit_latched), .B(steps_reg[0]), .C(\register_addr[1] ), 
         .Z(n30261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22851_3_lut.init = 16'hcaca;
    LUT4 i22853_3_lut (.A(Stepper_A_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22853_3_lut.init = 16'hcaca;
    LUT4 i22854_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22854_3_lut.init = 16'hcaca;
    LUT4 i14768_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14768_4_lut.init = 16'hc088;
    PFUMX i22852 (.BLUT(n30260), .ALUT(n30261), .C0(\register_addr[0] ), 
          .Z(n30262));
    PFUMX i22855 (.BLUT(n30263), .ALUT(n30264), .C0(\register_addr[1] ), 
          .Z(n30265));
    FD1P3AX int_step_182 (.D(n31917), .SP(n22_c), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i14769_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14769_4_lut.init = 16'hc088;
    LUT4 i14770_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14770_4_lut.init = 16'hc088;
    LUT4 i14771_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14771_4_lut.init = 16'hc088;
    LUT4 i22898_3_lut (.A(Stepper_A_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22898_3_lut.init = 16'hcaca;
    LUT4 i23177_4_lut (.A(n31911), .B(n32056), .C(n13323), .D(n32003), 
         .Z(n30489)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i23177_4_lut.init = 16'h0020;
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i22899_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22899_3_lut.init = 16'hcaca;
    LUT4 i14772_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14772_4_lut.init = 16'hc088;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_131), .C(n58_adj_132), .D(n50_adj_133), 
         .Z(n27766)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_134), .C(n54_adj_135), .D(n42_adj_136), 
         .Z(n62_adj_131)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i14773_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14773_4_lut.init = 16'hc088;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52_adj_137), .C(n38_adj_138), 
         .D(steps_reg[18]), .Z(n58_adj_132)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50_adj_133)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(steps_reg[9]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56_adj_139), .C(n46_adj_140), 
         .D(steps_reg[29]), .Z(n60_adj_134)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54_adj_135)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i14750_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14750_4_lut.init = 16'hc088;
    LUT4 i14751_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14751_4_lut.init = 16'hc088;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42_adj_136)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i14752_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14752_4_lut.init = 16'hc088;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(steps_reg[3]), .Z(n56_adj_139)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14753_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14753_4_lut.init = 16'hc088;
    LUT4 i14754_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14754_4_lut.init = 16'hc088;
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[6]), .Z(n46_adj_140)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i14755_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14755_4_lut.init = 16'hc088;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52_adj_137)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i14756_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14756_4_lut.init = 16'hc088;
    LUT4 i14757_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14757_4_lut.init = 16'hc088;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38_adj_138)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    PFUMX mux_1989_i4 (.BLUT(n8493[3]), .ALUT(n7348[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    LUT4 i14758_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14758_4_lut.init = 16'hc088;
    PFUMX mux_1989_i5 (.BLUT(n8493[4]), .ALUT(n7348[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    LUT4 i14759_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14759_4_lut.init = 16'hc088;
    PFUMX mux_1989_i6 (.BLUT(n8493[5]), .ALUT(n7348[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1989_i7 (.BLUT(n8493[6]), .ALUT(n7348[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    PFUMX mux_1989_i8 (.BLUT(n8494), .ALUT(n7348[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    ClockDivider_U9 step_clk_gen (.div_factor_reg({div_factor_reg}), .GND_net(GND_net), 
            .debug_c_c(debug_c_c), .n31903(n31903), .n16566(n16566), .step_clk(step_clk_c), 
            .n31991(n31991), .n8204(n8204), .n8238(n8238)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (div_factor_reg, GND_net, debug_c_c, n31903, 
            n16566, step_clk, n31991, n8204, n8238) /* synthesis syn_module_defined=1 */ ;
    input [31:0]div_factor_reg;
    input GND_net;
    input debug_c_c;
    input n31903;
    input n16566;
    output step_clk;
    input n31991;
    output n8204;
    output n8238;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27471, n27472, n27073;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n27074, n27072, n27071, n27470, n27469, n27468;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n26830, n27467, n27466, n27070, n27465, n27464, n27069, 
        n27463, n27068, n27462, n27461, n27460, n27067, n27066, 
        n27065, n27064, n27063, n27062, n8169;
    wire [31:0]n134;
    
    wire n26861, n26860, n26859, n26858, n26857, n26856, n26855, 
        n26854, n26853, n26852, n26851, n26850, n26849, n26848, 
        n26847, n26846, n26845, n26844, n26843, n26842, n26841, 
        n26840, n26839, n27320, n27319, n27318, n26838, n27317, 
        n27316, n27315, n27314, n27313, n26837, n26836, n27312, 
        n26835, n27311, n27310, n27309, n27308, n27307, n27306, 
        n27305, n26834, n26833, n26832, n27077, n27076, n26831, 
        n27075, n27475, n27474, n27473;
    
    CCU2D sub_2052_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27471), .COUT(n27472));
    defparam sub_2052_add_2_25.INIT0 = 16'hf555;
    defparam sub_2052_add_2_25.INIT1 = 16'hf555;
    defparam sub_2052_add_2_25.INJECT1_0 = "NO";
    defparam sub_2052_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27073), .COUT(n27074), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27072), .COUT(n27073), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27071), .COUT(n27072), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27470), .COUT(n27471));
    defparam sub_2052_add_2_23.INIT0 = 16'hf555;
    defparam sub_2052_add_2_23.INIT1 = 16'hf555;
    defparam sub_2052_add_2_23.INJECT1_0 = "NO";
    defparam sub_2052_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27469), .COUT(n27470));
    defparam sub_2052_add_2_21.INIT0 = 16'hf555;
    defparam sub_2052_add_2_21.INIT1 = 16'hf555;
    defparam sub_2052_add_2_21.INJECT1_0 = "NO";
    defparam sub_2052_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27468), .COUT(n27469));
    defparam sub_2052_add_2_19.INIT0 = 16'hf555;
    defparam sub_2052_add_2_19.INIT1 = 16'hf555;
    defparam sub_2052_add_2_19.INJECT1_0 = "NO";
    defparam sub_2052_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26830));
    defparam sub_2051_add_2_1.INIT0 = 16'h0000;
    defparam sub_2051_add_2_1.INIT1 = 16'h5999;
    defparam sub_2051_add_2_1.INJECT1_0 = "NO";
    defparam sub_2051_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27467), .COUT(n27468));
    defparam sub_2052_add_2_17.INIT0 = 16'hf555;
    defparam sub_2052_add_2_17.INIT1 = 16'hf555;
    defparam sub_2052_add_2_17.INJECT1_0 = "NO";
    defparam sub_2052_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27466), .COUT(n27467));
    defparam sub_2052_add_2_15.INIT0 = 16'hf555;
    defparam sub_2052_add_2_15.INIT1 = 16'hf555;
    defparam sub_2052_add_2_15.INJECT1_0 = "NO";
    defparam sub_2052_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27070), .COUT(n27071), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27465), .COUT(n27466));
    defparam sub_2052_add_2_13.INIT0 = 16'hf555;
    defparam sub_2052_add_2_13.INIT1 = 16'hf555;
    defparam sub_2052_add_2_13.INJECT1_0 = "NO";
    defparam sub_2052_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27464), .COUT(n27465));
    defparam sub_2052_add_2_11.INIT0 = 16'hf555;
    defparam sub_2052_add_2_11.INIT1 = 16'hf555;
    defparam sub_2052_add_2_11.INJECT1_0 = "NO";
    defparam sub_2052_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27069), .COUT(n27070), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27463), .COUT(n27464));
    defparam sub_2052_add_2_9.INIT0 = 16'hf555;
    defparam sub_2052_add_2_9.INIT1 = 16'hf555;
    defparam sub_2052_add_2_9.INJECT1_0 = "NO";
    defparam sub_2052_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27068), .COUT(n27069), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27462), .COUT(n27463));
    defparam sub_2052_add_2_7.INIT0 = 16'hf555;
    defparam sub_2052_add_2_7.INIT1 = 16'hf555;
    defparam sub_2052_add_2_7.INJECT1_0 = "NO";
    defparam sub_2052_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27461), .COUT(n27462));
    defparam sub_2052_add_2_5.INIT0 = 16'hf555;
    defparam sub_2052_add_2_5.INIT1 = 16'hf555;
    defparam sub_2052_add_2_5.INJECT1_0 = "NO";
    defparam sub_2052_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27460), .COUT(n27461));
    defparam sub_2052_add_2_3.INIT0 = 16'hf555;
    defparam sub_2052_add_2_3.INIT1 = 16'hf555;
    defparam sub_2052_add_2_3.INJECT1_0 = "NO";
    defparam sub_2052_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27460));
    defparam sub_2052_add_2_1.INIT0 = 16'h0000;
    defparam sub_2052_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2052_add_2_1.INJECT1_0 = "NO";
    defparam sub_2052_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27067), .COUT(n27068), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27066), .COUT(n27067), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27065), .COUT(n27066), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27064), .COUT(n27065), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27063), .COUT(n27064), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27062), .COUT(n27063), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27062), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8169), .CK(debug_c_c), .CD(n31991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2639__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i0.GSR = "ENABLED";
    CCU2D sub_2049_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26861), .S1(n8169));
    defparam sub_2049_add_2_33.INIT0 = 16'h5555;
    defparam sub_2049_add_2_33.INIT1 = 16'h0000;
    defparam sub_2049_add_2_33.INJECT1_0 = "NO";
    defparam sub_2049_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26860), .COUT(n26861));
    defparam sub_2049_add_2_31.INIT0 = 16'h5999;
    defparam sub_2049_add_2_31.INIT1 = 16'h5999;
    defparam sub_2049_add_2_31.INJECT1_0 = "NO";
    defparam sub_2049_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26859), .COUT(n26860));
    defparam sub_2049_add_2_29.INIT0 = 16'h5999;
    defparam sub_2049_add_2_29.INIT1 = 16'h5999;
    defparam sub_2049_add_2_29.INJECT1_0 = "NO";
    defparam sub_2049_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26858), .COUT(n26859));
    defparam sub_2049_add_2_27.INIT0 = 16'h5999;
    defparam sub_2049_add_2_27.INIT1 = 16'h5999;
    defparam sub_2049_add_2_27.INJECT1_0 = "NO";
    defparam sub_2049_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26857), .COUT(n26858));
    defparam sub_2049_add_2_25.INIT0 = 16'h5999;
    defparam sub_2049_add_2_25.INIT1 = 16'h5999;
    defparam sub_2049_add_2_25.INJECT1_0 = "NO";
    defparam sub_2049_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26856), .COUT(n26857));
    defparam sub_2049_add_2_23.INIT0 = 16'h5999;
    defparam sub_2049_add_2_23.INIT1 = 16'h5999;
    defparam sub_2049_add_2_23.INJECT1_0 = "NO";
    defparam sub_2049_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26855), .COUT(n26856));
    defparam sub_2049_add_2_21.INIT0 = 16'h5999;
    defparam sub_2049_add_2_21.INIT1 = 16'h5999;
    defparam sub_2049_add_2_21.INJECT1_0 = "NO";
    defparam sub_2049_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26854), .COUT(n26855));
    defparam sub_2049_add_2_19.INIT0 = 16'h5999;
    defparam sub_2049_add_2_19.INIT1 = 16'h5999;
    defparam sub_2049_add_2_19.INJECT1_0 = "NO";
    defparam sub_2049_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26853), .COUT(n26854));
    defparam sub_2049_add_2_17.INIT0 = 16'h5999;
    defparam sub_2049_add_2_17.INIT1 = 16'h5999;
    defparam sub_2049_add_2_17.INJECT1_0 = "NO";
    defparam sub_2049_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26852), .COUT(n26853));
    defparam sub_2049_add_2_15.INIT0 = 16'h5999;
    defparam sub_2049_add_2_15.INIT1 = 16'h5999;
    defparam sub_2049_add_2_15.INJECT1_0 = "NO";
    defparam sub_2049_add_2_15.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    CCU2D sub_2049_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26851), .COUT(n26852));
    defparam sub_2049_add_2_13.INIT0 = 16'h5999;
    defparam sub_2049_add_2_13.INIT1 = 16'h5999;
    defparam sub_2049_add_2_13.INJECT1_0 = "NO";
    defparam sub_2049_add_2_13.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31903), .CD(n16566), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31903), .PD(n16566), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2049_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26850), .COUT(n26851));
    defparam sub_2049_add_2_11.INIT0 = 16'h5999;
    defparam sub_2049_add_2_11.INIT1 = 16'h5999;
    defparam sub_2049_add_2_11.INJECT1_0 = "NO";
    defparam sub_2049_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26849), .COUT(n26850));
    defparam sub_2049_add_2_9.INIT0 = 16'h5999;
    defparam sub_2049_add_2_9.INIT1 = 16'h5999;
    defparam sub_2049_add_2_9.INJECT1_0 = "NO";
    defparam sub_2049_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26848), .COUT(n26849));
    defparam sub_2049_add_2_7.INIT0 = 16'h5999;
    defparam sub_2049_add_2_7.INIT1 = 16'h5999;
    defparam sub_2049_add_2_7.INJECT1_0 = "NO";
    defparam sub_2049_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26847), .COUT(n26848));
    defparam sub_2049_add_2_5.INIT0 = 16'h5999;
    defparam sub_2049_add_2_5.INIT1 = 16'h5999;
    defparam sub_2049_add_2_5.INJECT1_0 = "NO";
    defparam sub_2049_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26846), .COUT(n26847));
    defparam sub_2049_add_2_3.INIT0 = 16'h5999;
    defparam sub_2049_add_2_3.INIT1 = 16'h5999;
    defparam sub_2049_add_2_3.INJECT1_0 = "NO";
    defparam sub_2049_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2049_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26846));
    defparam sub_2049_add_2_1.INIT0 = 16'h0000;
    defparam sub_2049_add_2_1.INIT1 = 16'h5999;
    defparam sub_2049_add_2_1.INJECT1_0 = "NO";
    defparam sub_2049_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26845), .S1(n8204));
    defparam sub_2051_add_2_33.INIT0 = 16'h5999;
    defparam sub_2051_add_2_33.INIT1 = 16'h0000;
    defparam sub_2051_add_2_33.INJECT1_0 = "NO";
    defparam sub_2051_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26844), .COUT(n26845));
    defparam sub_2051_add_2_31.INIT0 = 16'h5999;
    defparam sub_2051_add_2_31.INIT1 = 16'h5999;
    defparam sub_2051_add_2_31.INJECT1_0 = "NO";
    defparam sub_2051_add_2_31.INJECT1_1 = "NO";
    FD1S3IX count_2639__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i1.GSR = "ENABLED";
    CCU2D sub_2051_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26843), .COUT(n26844));
    defparam sub_2051_add_2_29.INIT0 = 16'h5999;
    defparam sub_2051_add_2_29.INIT1 = 16'h5999;
    defparam sub_2051_add_2_29.INJECT1_0 = "NO";
    defparam sub_2051_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26842), .COUT(n26843));
    defparam sub_2051_add_2_27.INIT0 = 16'h5999;
    defparam sub_2051_add_2_27.INIT1 = 16'h5999;
    defparam sub_2051_add_2_27.INJECT1_0 = "NO";
    defparam sub_2051_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26841), .COUT(n26842));
    defparam sub_2051_add_2_25.INIT0 = 16'h5999;
    defparam sub_2051_add_2_25.INIT1 = 16'h5999;
    defparam sub_2051_add_2_25.INJECT1_0 = "NO";
    defparam sub_2051_add_2_25.INJECT1_1 = "NO";
    FD1S3IX count_2639__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i2.GSR = "ENABLED";
    FD1S3IX count_2639__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i3.GSR = "ENABLED";
    FD1S3IX count_2639__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i4.GSR = "ENABLED";
    FD1S3IX count_2639__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i5.GSR = "ENABLED";
    FD1S3IX count_2639__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i6.GSR = "ENABLED";
    FD1S3IX count_2639__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i7.GSR = "ENABLED";
    FD1S3IX count_2639__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i8.GSR = "ENABLED";
    FD1S3IX count_2639__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i9.GSR = "ENABLED";
    FD1S3IX count_2639__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i10.GSR = "ENABLED";
    FD1S3IX count_2639__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i11.GSR = "ENABLED";
    FD1S3IX count_2639__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i12.GSR = "ENABLED";
    FD1S3IX count_2639__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i13.GSR = "ENABLED";
    FD1S3IX count_2639__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i14.GSR = "ENABLED";
    FD1S3IX count_2639__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i15.GSR = "ENABLED";
    FD1S3IX count_2639__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i16.GSR = "ENABLED";
    FD1S3IX count_2639__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i17.GSR = "ENABLED";
    FD1S3IX count_2639__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i18.GSR = "ENABLED";
    FD1S3IX count_2639__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i19.GSR = "ENABLED";
    FD1S3IX count_2639__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i20.GSR = "ENABLED";
    FD1S3IX count_2639__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i21.GSR = "ENABLED";
    FD1S3IX count_2639__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i22.GSR = "ENABLED";
    FD1S3IX count_2639__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i23.GSR = "ENABLED";
    FD1S3IX count_2639__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i24.GSR = "ENABLED";
    FD1S3IX count_2639__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i25.GSR = "ENABLED";
    FD1S3IX count_2639__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i26.GSR = "ENABLED";
    FD1S3IX count_2639__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i27.GSR = "ENABLED";
    FD1S3IX count_2639__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i28.GSR = "ENABLED";
    FD1S3IX count_2639__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i29.GSR = "ENABLED";
    FD1S3IX count_2639__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i30.GSR = "ENABLED";
    FD1S3IX count_2639__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31903), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639__i31.GSR = "ENABLED";
    CCU2D sub_2051_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26840), .COUT(n26841));
    defparam sub_2051_add_2_23.INIT0 = 16'h5999;
    defparam sub_2051_add_2_23.INIT1 = 16'h5999;
    defparam sub_2051_add_2_23.INJECT1_0 = "NO";
    defparam sub_2051_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26839), .COUT(n26840));
    defparam sub_2051_add_2_21.INIT0 = 16'h5999;
    defparam sub_2051_add_2_21.INIT1 = 16'h5999;
    defparam sub_2051_add_2_21.INJECT1_0 = "NO";
    defparam sub_2051_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27320), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_33.INIT1 = 16'h0000;
    defparam count_2639_add_4_33.INJECT1_0 = "NO";
    defparam count_2639_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27319), .COUT(n27320), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_31.INJECT1_0 = "NO";
    defparam count_2639_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27318), .COUT(n27319), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_29.INJECT1_0 = "NO";
    defparam count_2639_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26838), .COUT(n26839));
    defparam sub_2051_add_2_19.INIT0 = 16'h5999;
    defparam sub_2051_add_2_19.INIT1 = 16'h5999;
    defparam sub_2051_add_2_19.INJECT1_0 = "NO";
    defparam sub_2051_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27317), .COUT(n27318), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_27.INJECT1_0 = "NO";
    defparam count_2639_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27316), .COUT(n27317), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_25.INJECT1_0 = "NO";
    defparam count_2639_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27315), .COUT(n27316), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_23.INJECT1_0 = "NO";
    defparam count_2639_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27314), .COUT(n27315), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_21.INJECT1_0 = "NO";
    defparam count_2639_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27313), .COUT(n27314), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_19.INJECT1_0 = "NO";
    defparam count_2639_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26837), .COUT(n26838));
    defparam sub_2051_add_2_17.INIT0 = 16'h5999;
    defparam sub_2051_add_2_17.INIT1 = 16'h5999;
    defparam sub_2051_add_2_17.INJECT1_0 = "NO";
    defparam sub_2051_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26836), .COUT(n26837));
    defparam sub_2051_add_2_15.INIT0 = 16'h5999;
    defparam sub_2051_add_2_15.INIT1 = 16'h5999;
    defparam sub_2051_add_2_15.INJECT1_0 = "NO";
    defparam sub_2051_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27312), .COUT(n27313), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_17.INJECT1_0 = "NO";
    defparam count_2639_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26835), .COUT(n26836));
    defparam sub_2051_add_2_13.INIT0 = 16'h5999;
    defparam sub_2051_add_2_13.INIT1 = 16'h5999;
    defparam sub_2051_add_2_13.INJECT1_0 = "NO";
    defparam sub_2051_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27311), .COUT(n27312), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_15.INJECT1_0 = "NO";
    defparam count_2639_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27310), .COUT(n27311), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_13.INJECT1_0 = "NO";
    defparam count_2639_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27309), .COUT(n27310), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_11.INJECT1_0 = "NO";
    defparam count_2639_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27308), .COUT(n27309), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_9.INJECT1_0 = "NO";
    defparam count_2639_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27307), .COUT(n27308), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_7.INJECT1_0 = "NO";
    defparam count_2639_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27306), .COUT(n27307), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_5.INJECT1_0 = "NO";
    defparam count_2639_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27305), .COUT(n27306), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2639_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2639_add_4_3.INJECT1_0 = "NO";
    defparam count_2639_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2639_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27305), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2639_add_4_1.INIT0 = 16'hF000;
    defparam count_2639_add_4_1.INIT1 = 16'h0555;
    defparam count_2639_add_4_1.INJECT1_0 = "NO";
    defparam count_2639_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26834), .COUT(n26835));
    defparam sub_2051_add_2_11.INIT0 = 16'h5999;
    defparam sub_2051_add_2_11.INIT1 = 16'h5999;
    defparam sub_2051_add_2_11.INJECT1_0 = "NO";
    defparam sub_2051_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26833), .COUT(n26834));
    defparam sub_2051_add_2_9.INIT0 = 16'h5999;
    defparam sub_2051_add_2_9.INIT1 = 16'h5999;
    defparam sub_2051_add_2_9.INJECT1_0 = "NO";
    defparam sub_2051_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26832), .COUT(n26833));
    defparam sub_2051_add_2_7.INIT0 = 16'h5999;
    defparam sub_2051_add_2_7.INIT1 = 16'h5999;
    defparam sub_2051_add_2_7.INJECT1_0 = "NO";
    defparam sub_2051_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27077), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27076), .COUT(n27077), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26831), .COUT(n26832));
    defparam sub_2051_add_2_5.INIT0 = 16'h5999;
    defparam sub_2051_add_2_5.INIT1 = 16'h5999;
    defparam sub_2051_add_2_5.INJECT1_0 = "NO";
    defparam sub_2051_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27075), .COUT(n27076), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2051_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26830), .COUT(n26831));
    defparam sub_2051_add_2_3.INIT0 = 16'h5999;
    defparam sub_2051_add_2_3.INIT1 = 16'h5999;
    defparam sub_2051_add_2_3.INJECT1_0 = "NO";
    defparam sub_2051_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27475), .S1(n8238));
    defparam sub_2052_add_2_33.INIT0 = 16'hf555;
    defparam sub_2052_add_2_33.INIT1 = 16'h0000;
    defparam sub_2052_add_2_33.INJECT1_0 = "NO";
    defparam sub_2052_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27474), .COUT(n27475));
    defparam sub_2052_add_2_31.INIT0 = 16'hf555;
    defparam sub_2052_add_2_31.INIT1 = 16'hf555;
    defparam sub_2052_add_2_31.INJECT1_0 = "NO";
    defparam sub_2052_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27473), .COUT(n27474));
    defparam sub_2052_add_2_29.INIT0 = 16'hf555;
    defparam sub_2052_add_2_29.INIT1 = 16'hf555;
    defparam sub_2052_add_2_29.INJECT1_0 = "NO";
    defparam sub_2052_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27472), .COUT(n27473));
    defparam sub_2052_add_2_27.INIT0 = 16'hf555;
    defparam sub_2052_add_2_27.INIT1 = 16'hf555;
    defparam sub_2052_add_2_27.INJECT1_0 = "NO";
    defparam sub_2052_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27074), .COUT(n27075), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (GND_net, clk_255kHz, debug_c_c, n241, n31991, 
            n7718, n30378, n14374, n30518, n27956, n30516, n27960, 
            n30381, n13735, n30505, n14315, n30445, n14358, n30514, 
            n27757, n2816, n7753, n30426, n14369, n30510, n27759, 
            n30520, n27883, n30512, n27758) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output clk_255kHz;
    input debug_c_c;
    input n241;
    input n31991;
    output n7718;
    input n30378;
    output n14374;
    input n30518;
    output n27956;
    input n30516;
    output n27960;
    input n30381;
    output n13735;
    input n30505;
    output n14315;
    input n30445;
    output n14358;
    input n30514;
    output n27757;
    input n2816;
    output n7753;
    input n30426;
    output n14369;
    input n30510;
    output n27759;
    input n30520;
    output n27883;
    input n30512;
    output n27758;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27267;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27268, n27266, n27265, n27264, n27263, n27262, n27261, 
        n27260, n27259, n27258, n27257, n27204, n27203, n27202, 
        n27201, n27200, n27199, n27198, n27197, n27196, n27195, 
        n27194, n27193, n27192, n27191, n27190, n27037, n27036, 
        n27035, n27034, n27033, n27032, n27031, n27030, n27029, 
        n27028, n27027, n27026, n27025, n27024, n27023, n27022, 
        n27272, n27271, n27270, n27269;
    
    CCU2D count_2633_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27267), .COUT(n27268), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_23.INJECT1_0 = "NO";
    defparam count_2633_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27266), .COUT(n27267), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_21.INJECT1_0 = "NO";
    defparam count_2633_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27265), .COUT(n27266), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_19.INJECT1_0 = "NO";
    defparam count_2633_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27264), .COUT(n27265), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_17.INJECT1_0 = "NO";
    defparam count_2633_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27263), .COUT(n27264), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_15.INJECT1_0 = "NO";
    defparam count_2633_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27262), .COUT(n27263), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_13.INJECT1_0 = "NO";
    defparam count_2633_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27261), .COUT(n27262), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_11.INJECT1_0 = "NO";
    defparam count_2633_add_4_11.INJECT1_1 = "NO";
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=544, LSE_RLINE=547 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D count_2633_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27260), .COUT(n27261), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_9.INJECT1_0 = "NO";
    defparam count_2633_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27259), .COUT(n27260), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_7.INJECT1_0 = "NO";
    defparam count_2633_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27258), .COUT(n27259), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_5.INJECT1_0 = "NO";
    defparam count_2633_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27257), .COUT(n27258), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_3.INJECT1_0 = "NO";
    defparam count_2633_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27257), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_1.INIT0 = 16'hF000;
    defparam count_2633_add_4_1.INIT1 = 16'h0555;
    defparam count_2633_add_4_1.INJECT1_0 = "NO";
    defparam count_2633_add_4_1.INJECT1_1 = "NO";
    LUT4 i23067_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30378), 
         .Z(n14374)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23067_2_lut_4_lut.init = 16'h1000;
    LUT4 i23207_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30518), 
         .Z(n27956)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23207_2_lut_4_lut.init = 16'h1000;
    LUT4 i23205_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30516), 
         .Z(n27960)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23205_2_lut_4_lut.init = 16'h1000;
    LUT4 i23070_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30381), 
         .Z(n13735)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23070_2_lut_4_lut.init = 16'h1000;
    LUT4 i23194_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30505), 
         .Z(n14315)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23194_2_lut_4_lut.init = 16'h1000;
    LUT4 i23134_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30445), 
         .Z(n14358)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23134_2_lut_4_lut.init = 16'h1000;
    LUT4 i23203_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30514), 
         .Z(n27757)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23203_2_lut_4_lut.init = 16'h1000;
    CCU2D add_20102_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27204), 
          .S1(n7718));
    defparam add_20102_32.INIT0 = 16'h5555;
    defparam add_20102_32.INIT1 = 16'h0000;
    defparam add_20102_32.INJECT1_0 = "NO";
    defparam add_20102_32.INJECT1_1 = "NO";
    CCU2D add_20102_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27203), .COUT(n27204));
    defparam add_20102_30.INIT0 = 16'h5555;
    defparam add_20102_30.INIT1 = 16'h5555;
    defparam add_20102_30.INJECT1_0 = "NO";
    defparam add_20102_30.INJECT1_1 = "NO";
    CCU2D add_20102_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27202), .COUT(n27203));
    defparam add_20102_28.INIT0 = 16'h5555;
    defparam add_20102_28.INIT1 = 16'h5555;
    defparam add_20102_28.INJECT1_0 = "NO";
    defparam add_20102_28.INJECT1_1 = "NO";
    CCU2D add_20102_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27201), .COUT(n27202));
    defparam add_20102_26.INIT0 = 16'h5555;
    defparam add_20102_26.INIT1 = 16'h5555;
    defparam add_20102_26.INJECT1_0 = "NO";
    defparam add_20102_26.INJECT1_1 = "NO";
    CCU2D add_20102_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27200), .COUT(n27201));
    defparam add_20102_24.INIT0 = 16'h5555;
    defparam add_20102_24.INIT1 = 16'h5555;
    defparam add_20102_24.INJECT1_0 = "NO";
    defparam add_20102_24.INJECT1_1 = "NO";
    CCU2D add_20102_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27199), .COUT(n27200));
    defparam add_20102_22.INIT0 = 16'h5555;
    defparam add_20102_22.INIT1 = 16'h5555;
    defparam add_20102_22.INJECT1_0 = "NO";
    defparam add_20102_22.INJECT1_1 = "NO";
    CCU2D add_20102_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27198), .COUT(n27199));
    defparam add_20102_20.INIT0 = 16'h5555;
    defparam add_20102_20.INIT1 = 16'h5555;
    defparam add_20102_20.INJECT1_0 = "NO";
    defparam add_20102_20.INJECT1_1 = "NO";
    CCU2D add_20102_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27197), .COUT(n27198));
    defparam add_20102_18.INIT0 = 16'h5555;
    defparam add_20102_18.INIT1 = 16'h5555;
    defparam add_20102_18.INJECT1_0 = "NO";
    defparam add_20102_18.INJECT1_1 = "NO";
    CCU2D add_20102_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27196), .COUT(n27197));
    defparam add_20102_16.INIT0 = 16'h5555;
    defparam add_20102_16.INIT1 = 16'h5555;
    defparam add_20102_16.INJECT1_0 = "NO";
    defparam add_20102_16.INJECT1_1 = "NO";
    CCU2D add_20102_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27195), .COUT(n27196));
    defparam add_20102_14.INIT0 = 16'h5555;
    defparam add_20102_14.INIT1 = 16'h5555;
    defparam add_20102_14.INJECT1_0 = "NO";
    defparam add_20102_14.INJECT1_1 = "NO";
    CCU2D add_20102_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27194), .COUT(n27195));
    defparam add_20102_12.INIT0 = 16'h5555;
    defparam add_20102_12.INIT1 = 16'h5555;
    defparam add_20102_12.INJECT1_0 = "NO";
    defparam add_20102_12.INJECT1_1 = "NO";
    CCU2D add_20102_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27193), .COUT(n27194));
    defparam add_20102_10.INIT0 = 16'h5555;
    defparam add_20102_10.INIT1 = 16'h5555;
    defparam add_20102_10.INJECT1_0 = "NO";
    defparam add_20102_10.INJECT1_1 = "NO";
    CCU2D add_20102_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27192), 
          .COUT(n27193));
    defparam add_20102_8.INIT0 = 16'h5555;
    defparam add_20102_8.INIT1 = 16'h5555;
    defparam add_20102_8.INJECT1_0 = "NO";
    defparam add_20102_8.INJECT1_1 = "NO";
    CCU2D add_20102_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27191), 
          .COUT(n27192));
    defparam add_20102_6.INIT0 = 16'h5555;
    defparam add_20102_6.INIT1 = 16'h5555;
    defparam add_20102_6.INJECT1_0 = "NO";
    defparam add_20102_6.INJECT1_1 = "NO";
    CCU2D add_20102_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27190), 
          .COUT(n27191));
    defparam add_20102_4.INIT0 = 16'h5555;
    defparam add_20102_4.INIT1 = 16'h5aaa;
    defparam add_20102_4.INJECT1_0 = "NO";
    defparam add_20102_4.INJECT1_1 = "NO";
    FD1S3IX count_2633__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2816), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i0.GSR = "ENABLED";
    CCU2D add_20102_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27190));
    defparam add_20102_2.INIT0 = 16'h7000;
    defparam add_20102_2.INIT1 = 16'h5aaa;
    defparam add_20102_2.INJECT1_0 = "NO";
    defparam add_20102_2.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27037), .S0(n7753));
    defparam sub_2029_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2029_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2029_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2029_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27036), .COUT(n27037));
    defparam sub_2029_add_2_32.INIT0 = 16'h5555;
    defparam sub_2029_add_2_32.INIT1 = 16'h5555;
    defparam sub_2029_add_2_32.INJECT1_0 = "NO";
    defparam sub_2029_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27035), .COUT(n27036));
    defparam sub_2029_add_2_30.INIT0 = 16'h5555;
    defparam sub_2029_add_2_30.INIT1 = 16'h5555;
    defparam sub_2029_add_2_30.INJECT1_0 = "NO";
    defparam sub_2029_add_2_30.INJECT1_1 = "NO";
    LUT4 i23115_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30426), 
         .Z(n14369)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23115_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_2029_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27034), .COUT(n27035));
    defparam sub_2029_add_2_28.INIT0 = 16'h5555;
    defparam sub_2029_add_2_28.INIT1 = 16'h5555;
    defparam sub_2029_add_2_28.INJECT1_0 = "NO";
    defparam sub_2029_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27033), .COUT(n27034));
    defparam sub_2029_add_2_26.INIT0 = 16'h5555;
    defparam sub_2029_add_2_26.INIT1 = 16'h5555;
    defparam sub_2029_add_2_26.INJECT1_0 = "NO";
    defparam sub_2029_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27032), .COUT(n27033));
    defparam sub_2029_add_2_24.INIT0 = 16'h5555;
    defparam sub_2029_add_2_24.INIT1 = 16'h5555;
    defparam sub_2029_add_2_24.INJECT1_0 = "NO";
    defparam sub_2029_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27031), .COUT(n27032));
    defparam sub_2029_add_2_22.INIT0 = 16'h5555;
    defparam sub_2029_add_2_22.INIT1 = 16'h5555;
    defparam sub_2029_add_2_22.INJECT1_0 = "NO";
    defparam sub_2029_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27030), .COUT(n27031));
    defparam sub_2029_add_2_20.INIT0 = 16'h5555;
    defparam sub_2029_add_2_20.INIT1 = 16'h5555;
    defparam sub_2029_add_2_20.INJECT1_0 = "NO";
    defparam sub_2029_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27029), .COUT(n27030));
    defparam sub_2029_add_2_18.INIT0 = 16'h5555;
    defparam sub_2029_add_2_18.INIT1 = 16'h5555;
    defparam sub_2029_add_2_18.INJECT1_0 = "NO";
    defparam sub_2029_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27028), .COUT(n27029));
    defparam sub_2029_add_2_16.INIT0 = 16'h5555;
    defparam sub_2029_add_2_16.INIT1 = 16'h5555;
    defparam sub_2029_add_2_16.INJECT1_0 = "NO";
    defparam sub_2029_add_2_16.INJECT1_1 = "NO";
    LUT4 i23199_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30510), 
         .Z(n27759)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23199_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_2029_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27027), .COUT(n27028));
    defparam sub_2029_add_2_14.INIT0 = 16'h5555;
    defparam sub_2029_add_2_14.INIT1 = 16'h5555;
    defparam sub_2029_add_2_14.INJECT1_0 = "NO";
    defparam sub_2029_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27026), .COUT(n27027));
    defparam sub_2029_add_2_12.INIT0 = 16'h5555;
    defparam sub_2029_add_2_12.INIT1 = 16'h5555;
    defparam sub_2029_add_2_12.INJECT1_0 = "NO";
    defparam sub_2029_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27025), .COUT(n27026));
    defparam sub_2029_add_2_10.INIT0 = 16'h5555;
    defparam sub_2029_add_2_10.INIT1 = 16'h5555;
    defparam sub_2029_add_2_10.INJECT1_0 = "NO";
    defparam sub_2029_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27024), .COUT(n27025));
    defparam sub_2029_add_2_8.INIT0 = 16'h5555;
    defparam sub_2029_add_2_8.INIT1 = 16'h5555;
    defparam sub_2029_add_2_8.INJECT1_0 = "NO";
    defparam sub_2029_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27023), .COUT(n27024));
    defparam sub_2029_add_2_6.INIT0 = 16'h5555;
    defparam sub_2029_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_2029_add_2_6.INJECT1_0 = "NO";
    defparam sub_2029_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27022), .COUT(n27023));
    defparam sub_2029_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2029_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_2029_add_2_4.INJECT1_0 = "NO";
    defparam sub_2029_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2029_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27022));
    defparam sub_2029_add_2_2.INIT0 = 16'h0000;
    defparam sub_2029_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2029_add_2_2.INJECT1_0 = "NO";
    defparam sub_2029_add_2_2.INJECT1_1 = "NO";
    LUT4 i23209_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30520), 
         .Z(n27883)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23209_2_lut_4_lut.init = 16'h1000;
    LUT4 i23201_2_lut_4_lut (.A(n31991), .B(clk_255kHz), .C(n7718), .D(n30512), 
         .Z(n27758)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23201_2_lut_4_lut.init = 16'h1000;
    FD1S3IX count_2633__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2816), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i1.GSR = "ENABLED";
    FD1S3IX count_2633__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2816), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i2.GSR = "ENABLED";
    FD1S3IX count_2633__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2816), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i3.GSR = "ENABLED";
    FD1S3IX count_2633__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2816), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i4.GSR = "ENABLED";
    FD1S3IX count_2633__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2816), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i5.GSR = "ENABLED";
    FD1S3IX count_2633__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2816), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i6.GSR = "ENABLED";
    FD1S3IX count_2633__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2816), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i7.GSR = "ENABLED";
    FD1S3IX count_2633__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2816), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i8.GSR = "ENABLED";
    FD1S3IX count_2633__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2816), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i9.GSR = "ENABLED";
    FD1S3IX count_2633__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i10.GSR = "ENABLED";
    FD1S3IX count_2633__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i11.GSR = "ENABLED";
    FD1S3IX count_2633__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i12.GSR = "ENABLED";
    FD1S3IX count_2633__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i13.GSR = "ENABLED";
    FD1S3IX count_2633__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i14.GSR = "ENABLED";
    FD1S3IX count_2633__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i15.GSR = "ENABLED";
    FD1S3IX count_2633__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i16.GSR = "ENABLED";
    FD1S3IX count_2633__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i17.GSR = "ENABLED";
    FD1S3IX count_2633__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i18.GSR = "ENABLED";
    FD1S3IX count_2633__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i19.GSR = "ENABLED";
    FD1S3IX count_2633__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i20.GSR = "ENABLED";
    FD1S3IX count_2633__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i21.GSR = "ENABLED";
    FD1S3IX count_2633__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i22.GSR = "ENABLED";
    FD1S3IX count_2633__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i23.GSR = "ENABLED";
    FD1S3IX count_2633__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i24.GSR = "ENABLED";
    FD1S3IX count_2633__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i25.GSR = "ENABLED";
    FD1S3IX count_2633__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i26.GSR = "ENABLED";
    FD1S3IX count_2633__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i27.GSR = "ENABLED";
    FD1S3IX count_2633__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i28.GSR = "ENABLED";
    FD1S3IX count_2633__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i29.GSR = "ENABLED";
    FD1S3IX count_2633__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i30.GSR = "ENABLED";
    FD1S3IX count_2633__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633__i31.GSR = "ENABLED";
    CCU2D count_2633_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27272), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_33.INIT1 = 16'h0000;
    defparam count_2633_add_4_33.INJECT1_0 = "NO";
    defparam count_2633_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27271), .COUT(n27272), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_31.INJECT1_0 = "NO";
    defparam count_2633_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27270), .COUT(n27271), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_29.INJECT1_0 = "NO";
    defparam count_2633_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27269), .COUT(n27270), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_27.INJECT1_0 = "NO";
    defparam count_2633_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2633_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27268), .COUT(n27269), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2633_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2633_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2633_add_4_25.INJECT1_0 = "NO";
    defparam count_2633_add_4_25.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ClockDividerP_SP(factor=120000) 
//

module \ClockDividerP_SP(factor=120000)  (debug_c_0, debug_c_c, n31991, 
            n2853, n30361, GND_net) /* synthesis syn_module_defined=1 */ ;
    output debug_c_0;
    input debug_c_c;
    input n31991;
    input n2853;
    output n30361;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(86[13:18])
    
    wire n21, n19, n20, n25, n36, n30, n38, n34, n26, n32, 
        n22, n28109;
    wire [31:0]n134;
    
    wire n31981, n30022, n30222, n30020, n30178, n30028, n27304, 
        n27303, n27302, n27301, n27300, n27299, n27298, n27297, 
        n27296, n27295, n27294, n27293, n27292, n27291, n27290, 
        n27289;
    
    LUT4 i9_4_lut (.A(count[5]), .B(count[16]), .C(count[12]), .D(count[14]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(count[7]), .B(count[15]), .C(count[4]), .D(count[10]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[1]), .B(count[0]), .C(count[2]), .D(count[3]), 
         .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[11]), .B(count[13]), .Z(n25)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(count[6]), .B(n36), .C(n30), .D(count[9]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(count[20]), .B(count[31]), .C(count[24]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(count[21]), .B(count[17]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i16_4_lut (.A(count[26]), .B(n32), .C(n22), .D(count[29]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(count[18]), .B(count[28]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(count[25]), .B(count[23]), .C(count[8]), .D(count[27]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[19]), .B(count[22]), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i2_2_lut.init = 16'heeee;
    FD1S3IX clk_o_13 (.D(n28109), .CK(debug_c_c), .CD(n31991), .Q(debug_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(88[9] 107[6])
    defparam clk_o_13.GSR = "ENABLED";
    FD1S3IX count_2634__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2853), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i0.GSR = "ENABLED";
    LUT4 i23122_4_lut_4_lut (.A(n31981), .B(n20), .C(n19), .D(n21), 
         .Z(n28109)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i23122_4_lut_4_lut.init = 16'h0001;
    LUT4 i23049_4_lut (.A(n31981), .B(n30022), .C(n30222), .D(n30020), 
         .Z(n30361)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i23049_4_lut.init = 16'h4000;
    LUT4 i22620_2_lut (.A(count[10]), .B(count[12]), .Z(n30022)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22620_2_lut.init = 16'h8888;
    LUT4 i22814_4_lut (.A(count[3]), .B(n30178), .C(n30028), .D(count[0]), 
         .Z(n30222)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22814_4_lut.init = 16'h8000;
    LUT4 i22618_2_lut (.A(count[2]), .B(count[5]), .Z(n30020)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22618_2_lut.init = 16'h8888;
    LUT4 i22770_4_lut (.A(count[1]), .B(count[16]), .C(count[4]), .D(count[15]), 
         .Z(n30178)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22770_4_lut.init = 16'h8000;
    LUT4 i22626_2_lut (.A(count[7]), .B(count[14]), .Z(n30028)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22626_2_lut.init = 16'h8888;
    FD1S3IX count_2634__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2853), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i1.GSR = "ENABLED";
    FD1S3IX count_2634__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2853), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i2.GSR = "ENABLED";
    FD1S3IX count_2634__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2853), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i3.GSR = "ENABLED";
    FD1S3IX count_2634__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2853), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i4.GSR = "ENABLED";
    FD1S3IX count_2634__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2853), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i5.GSR = "ENABLED";
    FD1S3IX count_2634__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2853), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i6.GSR = "ENABLED";
    FD1S3IX count_2634__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2853), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i7.GSR = "ENABLED";
    FD1S3IX count_2634__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2853), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i8.GSR = "ENABLED";
    FD1S3IX count_2634__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2853), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i9.GSR = "ENABLED";
    FD1S3IX count_2634__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i10.GSR = "ENABLED";
    FD1S3IX count_2634__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i11.GSR = "ENABLED";
    FD1S3IX count_2634__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i12.GSR = "ENABLED";
    FD1S3IX count_2634__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i13.GSR = "ENABLED";
    FD1S3IX count_2634__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i14.GSR = "ENABLED";
    FD1S3IX count_2634__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i15.GSR = "ENABLED";
    FD1S3IX count_2634__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i16.GSR = "ENABLED";
    FD1S3IX count_2634__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i17.GSR = "ENABLED";
    FD1S3IX count_2634__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i18.GSR = "ENABLED";
    FD1S3IX count_2634__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i19.GSR = "ENABLED";
    FD1S3IX count_2634__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i20.GSR = "ENABLED";
    FD1S3IX count_2634__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i21.GSR = "ENABLED";
    FD1S3IX count_2634__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i22.GSR = "ENABLED";
    FD1S3IX count_2634__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i23.GSR = "ENABLED";
    FD1S3IX count_2634__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i24.GSR = "ENABLED";
    FD1S3IX count_2634__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i25.GSR = "ENABLED";
    FD1S3IX count_2634__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i26.GSR = "ENABLED";
    FD1S3IX count_2634__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i27.GSR = "ENABLED";
    FD1S3IX count_2634__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i28.GSR = "ENABLED";
    FD1S3IX count_2634__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i29.GSR = "ENABLED";
    FD1S3IX count_2634__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i30.GSR = "ENABLED";
    FD1S3IX count_2634__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2853), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634__i31.GSR = "ENABLED";
    CCU2D count_2634_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27304), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_33.INIT1 = 16'h0000;
    defparam count_2634_add_4_33.INJECT1_0 = "NO";
    defparam count_2634_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27303), .COUT(n27304), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_31.INJECT1_0 = "NO";
    defparam count_2634_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27302), .COUT(n27303), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_29.INJECT1_0 = "NO";
    defparam count_2634_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27301), .COUT(n27302), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_27.INJECT1_0 = "NO";
    defparam count_2634_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27300), .COUT(n27301), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_25.INJECT1_0 = "NO";
    defparam count_2634_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27299), .COUT(n27300), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_23.INJECT1_0 = "NO";
    defparam count_2634_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27298), .COUT(n27299), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_21.INJECT1_0 = "NO";
    defparam count_2634_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27297), .COUT(n27298), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_19.INJECT1_0 = "NO";
    defparam count_2634_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27296), .COUT(n27297), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_17.INJECT1_0 = "NO";
    defparam count_2634_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27295), .COUT(n27296), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_15.INJECT1_0 = "NO";
    defparam count_2634_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27294), .COUT(n27295), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_13.INJECT1_0 = "NO";
    defparam count_2634_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27293), .COUT(n27294), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_11.INJECT1_0 = "NO";
    defparam count_2634_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27292), .COUT(n27293), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_9.INJECT1_0 = "NO";
    defparam count_2634_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27291), .COUT(n27292), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_7.INJECT1_0 = "NO";
    defparam count_2634_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27290), .COUT(n27291), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_5.INJECT1_0 = "NO";
    defparam count_2634_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27289), .COUT(n27290), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2634_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2634_add_4_3.INJECT1_0 = "NO";
    defparam count_2634_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2634_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27289), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2634_add_4_1.INIT0 = 16'hF000;
    defparam count_2634_add_4_1.INIT1 = 16'h0555;
    defparam count_2634_add_4_1.INJECT1_0 = "NO";
    defparam count_2634_add_4_1.INJECT1_1 = "NO";
    LUT4 i19_4_lut_rep_364 (.A(n25), .B(n38), .C(n34), .D(n26), .Z(n31981)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i19_4_lut_rep_364.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (read_value, debug_c_c, n13876, 
            GND_net, VCC_net, Stepper_Z_nFault_c, \read_size[0] , n29175, 
            n31991, Stepper_Z_M0_c_0, n110, n579, prev_step_clk, step_clk, 
            limit_latched, prev_limit_latched, n13698, prev_select, 
            n31982, databus, n3984, \register_addr[1] , \register_addr[0] , 
            n27787, \read_size[2] , n29174, Stepper_Z_M1_c_1, n13693, 
            Stepper_Z_M2_c_2, Stepper_Z_Dir_c, Stepper_Z_En_c, \control_reg[7] , 
            n11020, n9139, n32, n22, n31918, limit_c_2, Stepper_Z_Step_c, 
            n8485, n8100, n31902, n16565, n8134) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n13876;
    input GND_net;
    input VCC_net;
    input Stepper_Z_nFault_c;
    output \read_size[0] ;
    input n29175;
    input n31991;
    output Stepper_Z_M0_c_0;
    input n110;
    input n579;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    input n13698;
    output prev_select;
    input n31982;
    input [31:0]databus;
    input n3984;
    input \register_addr[1] ;
    input \register_addr[0] ;
    output n27787;
    output \read_size[2] ;
    input n29174;
    output Stepper_Z_M1_c_1;
    input n13693;
    output Stepper_Z_M2_c_2;
    output Stepper_Z_Dir_c;
    output Stepper_Z_En_c;
    output \control_reg[7] ;
    input n11020;
    input n9139;
    input n32;
    input n22;
    input n31918;
    input limit_c_2;
    output Stepper_Z_Step_c;
    input n8485;
    output n8100;
    input n31902;
    input n16565;
    output n8134;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n30343, fault_latched;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n3985;
    
    wire n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]n224;
    wire [31:0]n100;
    
    wire n30341, n30342, n30304, n30301, n49, n62, n58, n50;
    wire [31:0]n99;
    
    wire n16, n30302, n30303;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n27157, n27156, n27155, n41, n60, n54, n42_adj_117, n52, 
        n38_adj_118, n27154, n27153, n27152, n27151, n27150, n27149, 
        n27148, n27147, n27146, n27145, n27144, n27143, n27142, 
        n56, n46_adj_119, n23, int_step, n30299, n30300;
    wire [7:0]n8484;
    wire [31:0]n7034;
    
    FD1P3IX read_value__i0 (.D(n30343), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n29175), .SP(n13876), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3985[0]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n110), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13698), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31982), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3985[31]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3985[30]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3985[29]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3985[28]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3985[27]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3985[26]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3985[25]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3985[24]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3985[23]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3985[22]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3985[21]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    LUT4 mux_1559_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3984), .Z(n3985[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i8_3_lut.init = 16'hcaca;
    LUT4 i14778_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14778_4_lut.init = 16'hc088;
    LUT4 i14779_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14779_4_lut.init = 16'hc088;
    LUT4 i14780_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14780_4_lut.init = 16'hc088;
    LUT4 i14781_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14781_4_lut.init = 16'hc088;
    LUT4 i14782_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14782_4_lut.init = 16'hc088;
    LUT4 i14783_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14783_4_lut.init = 16'hc088;
    LUT4 i14784_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14784_4_lut.init = 16'hc088;
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[24]), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i14785_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14785_4_lut.init = 16'hc088;
    LUT4 i14786_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14786_4_lut.init = 16'hc088;
    LUT4 i14787_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14787_4_lut.init = 16'hc088;
    LUT4 i14788_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14788_4_lut.init = 16'hc088;
    LUT4 i14789_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14789_4_lut.init = 16'hc088;
    LUT4 i14790_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14790_4_lut.init = 16'hc088;
    LUT4 i14791_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14791_4_lut.init = 16'hc088;
    LUT4 i22931_3_lut (.A(Stepper_Z_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22931_3_lut.init = 16'hcaca;
    LUT4 i22932_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22932_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n13876), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30304), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30301), .SP(n13876), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1559_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3984), .Z(n3985[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i7_3_lut.init = 16'hcaca;
    PFUMX i22933 (.BLUT(n30341), .ALUT(n30342), .C0(\register_addr[1] ), 
          .Z(n30343));
    LUT4 mux_1559_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3984), .Z(n3985[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3984), .Z(n3985[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i5_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27787)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 mux_1559_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3984), .Z(n3985[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i4_3_lut.init = 16'hcaca;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[8]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    FD1P3AX read_value__i15 (.D(n99[15]), .SP(n13876), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_237 (.A(\register_addr[1] ), .B(div_factor_reg[16]), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n16)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_237.init = 16'ha088;
    LUT4 i15325_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n99[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i15325_4_lut.init = 16'hc088;
    FD1S3IX steps_reg__i20 (.D(n3985[20]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3985[19]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3985[18]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3985[17]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3985[16]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3985[15]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3985[14]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3985[13]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3985[12]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3985[11]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3985[10]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3985[9]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3985[8]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3985[7]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3985[6]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3985[5]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3985[4]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3985[3]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3985[2]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3985[1]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n29174), .SP(n13876), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i15324_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n99[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i15324_4_lut.init = 16'hc088;
    LUT4 mux_1559_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3984), .Z(n3985[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i3_3_lut.init = 16'hcaca;
    PFUMX i22894 (.BLUT(n30302), .ALUT(n30303), .C0(\register_addr[0] ), 
          .Z(n30304));
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13693), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13693), .CD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13693), .PD(n31991), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13693), .CD(n31991), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13693), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13693), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13693), .CD(n11020), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9139), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9139), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9139), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9139), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9139), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9139), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9139), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9139), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i15326_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n99[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i15326_4_lut.init = 16'hc088;
    LUT4 mux_1559_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3984), 
         .Z(n3985[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3984), 
         .Z(n3985[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3984), 
         .Z(n3985[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3984), 
         .Z(n3985[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3984), 
         .Z(n3985[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3984), 
         .Z(n3985[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3984), 
         .Z(n3985[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3984), 
         .Z(n3985[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3984), 
         .Z(n3985[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3984), .Z(n3985[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3984), .Z(n3985[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3984), 
         .Z(n3985[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3984), 
         .Z(n3985[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i11_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27157), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    LUT4 mux_1559_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3984), .Z(n3985[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i10_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27156), .COUT(n27157), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27155), .COUT(n27156), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42_adj_117), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38_adj_118), .D(steps_reg[16]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 mux_1559_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3984), 
         .Z(n3985[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i23_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27154), .COUT(n27155), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27153), .COUT(n27154), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27152), .COUT(n27153), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27151), .COUT(n27152), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27150), .COUT(n27151), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27149), .COUT(n27150), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27148), .COUT(n27149), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27147), .COUT(n27148), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    LUT4 mux_1559_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3984), 
         .Z(n3985[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i22_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27146), .COUT(n27147), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27145), .COUT(n27146), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27144), .COUT(n27145), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27143), .COUT(n27144), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27142), .COUT(n27143), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27142), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[18]), .B(steps_reg[0]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[12]), .B(n56), .C(n46_adj_119), .D(steps_reg[17]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[29]), .B(steps_reg[4]), .C(steps_reg[24]), 
         .D(steps_reg[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i15323_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n99[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i15323_4_lut.init = 16'hc088;
    LUT4 i10_2_lut (.A(steps_reg[25]), .B(steps_reg[26]), .Z(n42_adj_117)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[5]), .B(steps_reg[10]), .C(steps_reg[6]), 
         .D(steps_reg[3]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_238 (.A(div_factor_reg[20]), .B(\register_addr[1] ), 
         .C(steps_reg[20]), .D(\register_addr[0] ), .Z(n23)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    defparam i1_4_lut_adj_238.init = 16'hc088;
    LUT4 i14_2_lut (.A(steps_reg[22]), .B(steps_reg[2]), .Z(n46_adj_119)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[28]), .B(steps_reg[7]), .C(steps_reg[30]), 
         .D(steps_reg[20]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[1]), .B(steps_reg[13]), .Z(n38_adj_118)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    FD1P3AX read_value__i16 (.D(n16), .SP(n13876), .CK(debug_c_c), .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n99[17]), .SP(n13876), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n99[18]), .SP(n13876), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    LUT4 i15322_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n99[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i15322_4_lut.init = 16'hc088;
    FD1P3AX read_value__i19 (.D(n99[19]), .SP(n13876), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n23), .SP(n13876), .CK(debug_c_c), .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n99[21]), .SP(n13876), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    LUT4 i15321_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n99[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i15321_4_lut.init = 16'hc088;
    LUT4 i15320_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n99[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i15320_4_lut.init = 16'hc088;
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n99[22]), .SP(n13876), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n13698), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n99[23]), .SP(n13876), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=614, LSE_RLINE=627 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n31918), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1559_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3984), .Z(n3985[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i1_3_lut.init = 16'hcaca;
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    PFUMX i22891 (.BLUT(n30299), .ALUT(n30300), .C0(\register_addr[0] ), 
          .Z(n30301));
    PFUMX mux_1963_i4 (.BLUT(n8484[3]), .ALUT(n7034[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    LUT4 i22889_3_lut (.A(Stepper_Z_M1_c_1), .B(div_factor_reg[1]), .C(\register_addr[1] ), 
         .Z(n30299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22889_3_lut.init = 16'hcaca;
    LUT4 i22890_3_lut (.A(fault_latched), .B(steps_reg[1]), .C(\register_addr[1] ), 
         .Z(n30300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22890_3_lut.init = 16'hcaca;
    PFUMX mux_1963_i5 (.BLUT(n8484[4]), .ALUT(n7034[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1963_i6 (.BLUT(n8484[5]), .ALUT(n7034[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1963_i7 (.BLUT(n8484[6]), .ALUT(n7034[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i14777_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8484[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14777_2_lut.init = 16'h2222;
    LUT4 mux_1959_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7034[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1959_i4_3_lut.init = 16'hcaca;
    LUT4 i14776_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8484[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14776_2_lut.init = 16'h2222;
    LUT4 mux_1959_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7034[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1959_i5_3_lut.init = 16'hcaca;
    LUT4 i14775_2_lut (.A(Stepper_Z_Dir_c), .B(\register_addr[0] ), .Z(n8484[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14775_2_lut.init = 16'h2222;
    LUT4 mux_1959_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7034[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1959_i6_3_lut.init = 16'hcaca;
    PFUMX mux_1963_i8 (.BLUT(n8485), .ALUT(n7034[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    LUT4 i14774_2_lut (.A(Stepper_Z_En_c), .B(\register_addr[0] ), .Z(n8484[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14774_2_lut.init = 16'h2222;
    LUT4 mux_1959_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7034[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1959_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3984), 
         .Z(n3985[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1959_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n7034[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1959_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3984), 
         .Z(n3985[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3984), 
         .Z(n3985[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3984), 
         .Z(n3985[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3984), 
         .Z(n3985[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3984), 
         .Z(n3985[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3984), 
         .Z(n3985[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3984), 
         .Z(n3985[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3984), 
         .Z(n3985[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1559_i24_3_lut.init = 16'hcaca;
    LUT4 i22892_3_lut (.A(Stepper_Z_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22892_3_lut.init = 16'hcaca;
    LUT4 i22893_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22893_3_lut.init = 16'hcaca;
    ClockDivider step_clk_gen (.GND_net(GND_net), .n8100(n8100), .debug_c_c(debug_c_c), 
            .n31902(n31902), .n16565(n16565), .div_factor_reg({div_factor_reg}), 
            .step_clk(step_clk), .n31991(n31991), .n8134(n8134)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (GND_net, n8100, debug_c_c, n31902, n16565, div_factor_reg, 
            step_clk, n31991, n8134) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n8100;
    input debug_c_c;
    input n31902;
    input n16565;
    input [31:0]div_factor_reg;
    output step_clk;
    input n31991;
    output n8134;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26898;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26899, n26897, n26896, n26895, n26894, n26893;
    wire [31:0]n40;
    
    wire n26892, n26891, n26890, n26889, n26888, n8065, n26887, 
        n26886, n26885, n26884, n26883, n26882, n26881, n26880, 
        n26879, n26878, n26877, n26876, n26875, n26874, n26873;
    wire [31:0]n134;
    
    wire n26872, n26871, n26870, n26869, n26868, n26867, n26866, 
        n26865, n26864, n26863, n26862, n27093, n27092, n27091, 
        n27090, n27089, n27088, n26909, n27087, n27288, n27287, 
        n27286, n26908, n26907, n27285, n27086, n27284, n27085, 
        n26906, n27084, n27083, n26905, n27283, n27082, n26904, 
        n27282, n27281, n26903, n27081, n27280, n27080, n27079, 
        n27078, n27279, n27278, n27277, n27276, n27275, n27274, 
        n27273, n26902, n26901, n26900;
    
    CCU2D sub_2044_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26898), .COUT(n26899));
    defparam sub_2044_add_2_11.INIT0 = 16'h5999;
    defparam sub_2044_add_2_11.INIT1 = 16'h5999;
    defparam sub_2044_add_2_11.INJECT1_0 = "NO";
    defparam sub_2044_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26897), .COUT(n26898));
    defparam sub_2044_add_2_9.INIT0 = 16'h5999;
    defparam sub_2044_add_2_9.INIT1 = 16'h5999;
    defparam sub_2044_add_2_9.INJECT1_0 = "NO";
    defparam sub_2044_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26896), .COUT(n26897));
    defparam sub_2044_add_2_7.INIT0 = 16'h5999;
    defparam sub_2044_add_2_7.INIT1 = 16'h5999;
    defparam sub_2044_add_2_7.INJECT1_0 = "NO";
    defparam sub_2044_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26895), .COUT(n26896));
    defparam sub_2044_add_2_5.INIT0 = 16'h5999;
    defparam sub_2044_add_2_5.INIT1 = 16'h5999;
    defparam sub_2044_add_2_5.INJECT1_0 = "NO";
    defparam sub_2044_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26894), .COUT(n26895));
    defparam sub_2044_add_2_3.INIT0 = 16'h5999;
    defparam sub_2044_add_2_3.INIT1 = 16'h5999;
    defparam sub_2044_add_2_3.INJECT1_0 = "NO";
    defparam sub_2044_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26894));
    defparam sub_2044_add_2_1.INIT0 = 16'h0000;
    defparam sub_2044_add_2_1.INIT1 = 16'h5999;
    defparam sub_2044_add_2_1.INJECT1_0 = "NO";
    defparam sub_2044_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26893), .S1(n8100));
    defparam sub_2046_add_2_33.INIT0 = 16'h5999;
    defparam sub_2046_add_2_33.INIT1 = 16'h0000;
    defparam sub_2046_add_2_33.INJECT1_0 = "NO";
    defparam sub_2046_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26892), .COUT(n26893));
    defparam sub_2046_add_2_31.INIT0 = 16'h5999;
    defparam sub_2046_add_2_31.INIT1 = 16'h5999;
    defparam sub_2046_add_2_31.INJECT1_0 = "NO";
    defparam sub_2046_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26891), .COUT(n26892));
    defparam sub_2046_add_2_29.INIT0 = 16'h5999;
    defparam sub_2046_add_2_29.INIT1 = 16'h5999;
    defparam sub_2046_add_2_29.INJECT1_0 = "NO";
    defparam sub_2046_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26890), .COUT(n26891));
    defparam sub_2046_add_2_27.INIT0 = 16'h5999;
    defparam sub_2046_add_2_27.INIT1 = 16'h5999;
    defparam sub_2046_add_2_27.INJECT1_0 = "NO";
    defparam sub_2046_add_2_27.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2046_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26889), .COUT(n26890));
    defparam sub_2046_add_2_25.INIT0 = 16'h5999;
    defparam sub_2046_add_2_25.INIT1 = 16'h5999;
    defparam sub_2046_add_2_25.INJECT1_0 = "NO";
    defparam sub_2046_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26888), .COUT(n26889));
    defparam sub_2046_add_2_23.INIT0 = 16'h5999;
    defparam sub_2046_add_2_23.INIT1 = 16'h5999;
    defparam sub_2046_add_2_23.INJECT1_0 = "NO";
    defparam sub_2046_add_2_23.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8065), .CK(debug_c_c), .CD(n31991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2046_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26887), .COUT(n26888));
    defparam sub_2046_add_2_21.INIT0 = 16'h5999;
    defparam sub_2046_add_2_21.INIT1 = 16'h5999;
    defparam sub_2046_add_2_21.INJECT1_0 = "NO";
    defparam sub_2046_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26886), .COUT(n26887));
    defparam sub_2046_add_2_19.INIT0 = 16'h5999;
    defparam sub_2046_add_2_19.INIT1 = 16'h5999;
    defparam sub_2046_add_2_19.INJECT1_0 = "NO";
    defparam sub_2046_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26885), .COUT(n26886));
    defparam sub_2046_add_2_17.INIT0 = 16'h5999;
    defparam sub_2046_add_2_17.INIT1 = 16'h5999;
    defparam sub_2046_add_2_17.INJECT1_0 = "NO";
    defparam sub_2046_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26884), .COUT(n26885));
    defparam sub_2046_add_2_15.INIT0 = 16'h5999;
    defparam sub_2046_add_2_15.INIT1 = 16'h5999;
    defparam sub_2046_add_2_15.INJECT1_0 = "NO";
    defparam sub_2046_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26883), .COUT(n26884));
    defparam sub_2046_add_2_13.INIT0 = 16'h5999;
    defparam sub_2046_add_2_13.INIT1 = 16'h5999;
    defparam sub_2046_add_2_13.INJECT1_0 = "NO";
    defparam sub_2046_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26882), .COUT(n26883));
    defparam sub_2046_add_2_11.INIT0 = 16'h5999;
    defparam sub_2046_add_2_11.INIT1 = 16'h5999;
    defparam sub_2046_add_2_11.INJECT1_0 = "NO";
    defparam sub_2046_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26881), .COUT(n26882));
    defparam sub_2046_add_2_9.INIT0 = 16'h5999;
    defparam sub_2046_add_2_9.INIT1 = 16'h5999;
    defparam sub_2046_add_2_9.INJECT1_0 = "NO";
    defparam sub_2046_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26880), .COUT(n26881));
    defparam sub_2046_add_2_7.INIT0 = 16'h5999;
    defparam sub_2046_add_2_7.INIT1 = 16'h5999;
    defparam sub_2046_add_2_7.INJECT1_0 = "NO";
    defparam sub_2046_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26879), .COUT(n26880));
    defparam sub_2046_add_2_5.INIT0 = 16'h5999;
    defparam sub_2046_add_2_5.INIT1 = 16'h5999;
    defparam sub_2046_add_2_5.INJECT1_0 = "NO";
    defparam sub_2046_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26878), .COUT(n26879));
    defparam sub_2046_add_2_3.INIT0 = 16'h5999;
    defparam sub_2046_add_2_3.INIT1 = 16'h5999;
    defparam sub_2046_add_2_3.INJECT1_0 = "NO";
    defparam sub_2046_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2046_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26878));
    defparam sub_2046_add_2_1.INIT0 = 16'h0000;
    defparam sub_2046_add_2_1.INIT1 = 16'h5999;
    defparam sub_2046_add_2_1.INJECT1_0 = "NO";
    defparam sub_2046_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26877), .S1(n8134));
    defparam sub_2047_add_2_33.INIT0 = 16'hf555;
    defparam sub_2047_add_2_33.INIT1 = 16'h0000;
    defparam sub_2047_add_2_33.INJECT1_0 = "NO";
    defparam sub_2047_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26876), .COUT(n26877));
    defparam sub_2047_add_2_31.INIT0 = 16'hf555;
    defparam sub_2047_add_2_31.INIT1 = 16'hf555;
    defparam sub_2047_add_2_31.INJECT1_0 = "NO";
    defparam sub_2047_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26875), .COUT(n26876));
    defparam sub_2047_add_2_29.INIT0 = 16'hf555;
    defparam sub_2047_add_2_29.INIT1 = 16'hf555;
    defparam sub_2047_add_2_29.INJECT1_0 = "NO";
    defparam sub_2047_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26874), .COUT(n26875));
    defparam sub_2047_add_2_27.INIT0 = 16'hf555;
    defparam sub_2047_add_2_27.INIT1 = 16'hf555;
    defparam sub_2047_add_2_27.INJECT1_0 = "NO";
    defparam sub_2047_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26873), .COUT(n26874));
    defparam sub_2047_add_2_25.INIT0 = 16'hf555;
    defparam sub_2047_add_2_25.INIT1 = 16'hf555;
    defparam sub_2047_add_2_25.INJECT1_0 = "NO";
    defparam sub_2047_add_2_25.INJECT1_1 = "NO";
    FD1S3IX count_2638__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i0.GSR = "ENABLED";
    CCU2D sub_2047_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26872), .COUT(n26873));
    defparam sub_2047_add_2_23.INIT0 = 16'hf555;
    defparam sub_2047_add_2_23.INIT1 = 16'hf555;
    defparam sub_2047_add_2_23.INJECT1_0 = "NO";
    defparam sub_2047_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26871), .COUT(n26872));
    defparam sub_2047_add_2_21.INIT0 = 16'hf555;
    defparam sub_2047_add_2_21.INIT1 = 16'hf555;
    defparam sub_2047_add_2_21.INJECT1_0 = "NO";
    defparam sub_2047_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26870), .COUT(n26871));
    defparam sub_2047_add_2_19.INIT0 = 16'hf555;
    defparam sub_2047_add_2_19.INIT1 = 16'hf555;
    defparam sub_2047_add_2_19.INJECT1_0 = "NO";
    defparam sub_2047_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26869), .COUT(n26870));
    defparam sub_2047_add_2_17.INIT0 = 16'hf555;
    defparam sub_2047_add_2_17.INIT1 = 16'hf555;
    defparam sub_2047_add_2_17.INJECT1_0 = "NO";
    defparam sub_2047_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26868), .COUT(n26869));
    defparam sub_2047_add_2_15.INIT0 = 16'hf555;
    defparam sub_2047_add_2_15.INIT1 = 16'hf555;
    defparam sub_2047_add_2_15.INJECT1_0 = "NO";
    defparam sub_2047_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26867), .COUT(n26868));
    defparam sub_2047_add_2_13.INIT0 = 16'hf555;
    defparam sub_2047_add_2_13.INIT1 = 16'hf555;
    defparam sub_2047_add_2_13.INJECT1_0 = "NO";
    defparam sub_2047_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26866), .COUT(n26867));
    defparam sub_2047_add_2_11.INIT0 = 16'hf555;
    defparam sub_2047_add_2_11.INIT1 = 16'hf555;
    defparam sub_2047_add_2_11.INJECT1_0 = "NO";
    defparam sub_2047_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26865), .COUT(n26866));
    defparam sub_2047_add_2_9.INIT0 = 16'hf555;
    defparam sub_2047_add_2_9.INIT1 = 16'hf555;
    defparam sub_2047_add_2_9.INJECT1_0 = "NO";
    defparam sub_2047_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26864), .COUT(n26865));
    defparam sub_2047_add_2_7.INIT0 = 16'hf555;
    defparam sub_2047_add_2_7.INIT1 = 16'hf555;
    defparam sub_2047_add_2_7.INJECT1_0 = "NO";
    defparam sub_2047_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26863), .COUT(n26864));
    defparam sub_2047_add_2_5.INIT0 = 16'hf555;
    defparam sub_2047_add_2_5.INIT1 = 16'hf555;
    defparam sub_2047_add_2_5.INJECT1_0 = "NO";
    defparam sub_2047_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26862), .COUT(n26863));
    defparam sub_2047_add_2_3.INIT0 = 16'hf555;
    defparam sub_2047_add_2_3.INIT1 = 16'hf555;
    defparam sub_2047_add_2_3.INJECT1_0 = "NO";
    defparam sub_2047_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26862));
    defparam sub_2047_add_2_1.INIT0 = 16'h0000;
    defparam sub_2047_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2047_add_2_1.INJECT1_0 = "NO";
    defparam sub_2047_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31902), .CD(n16565), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31902), .PD(n16565), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1S3IX count_2638__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i1.GSR = "ENABLED";
    FD1S3IX count_2638__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i2.GSR = "ENABLED";
    FD1S3IX count_2638__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i3.GSR = "ENABLED";
    FD1S3IX count_2638__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i4.GSR = "ENABLED";
    FD1S3IX count_2638__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i5.GSR = "ENABLED";
    FD1S3IX count_2638__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i6.GSR = "ENABLED";
    FD1S3IX count_2638__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i7.GSR = "ENABLED";
    FD1S3IX count_2638__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i8.GSR = "ENABLED";
    FD1S3IX count_2638__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i9.GSR = "ENABLED";
    FD1S3IX count_2638__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i10.GSR = "ENABLED";
    FD1S3IX count_2638__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i11.GSR = "ENABLED";
    FD1S3IX count_2638__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i12.GSR = "ENABLED";
    FD1S3IX count_2638__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i13.GSR = "ENABLED";
    FD1S3IX count_2638__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i14.GSR = "ENABLED";
    FD1S3IX count_2638__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i15.GSR = "ENABLED";
    FD1S3IX count_2638__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i16.GSR = "ENABLED";
    FD1S3IX count_2638__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i17.GSR = "ENABLED";
    FD1S3IX count_2638__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i18.GSR = "ENABLED";
    FD1S3IX count_2638__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i19.GSR = "ENABLED";
    FD1S3IX count_2638__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i20.GSR = "ENABLED";
    FD1S3IX count_2638__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i21.GSR = "ENABLED";
    FD1S3IX count_2638__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i22.GSR = "ENABLED";
    FD1S3IX count_2638__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i23.GSR = "ENABLED";
    FD1S3IX count_2638__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i24.GSR = "ENABLED";
    FD1S3IX count_2638__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i25.GSR = "ENABLED";
    FD1S3IX count_2638__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i26.GSR = "ENABLED";
    FD1S3IX count_2638__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i27.GSR = "ENABLED";
    FD1S3IX count_2638__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i28.GSR = "ENABLED";
    FD1S3IX count_2638__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i29.GSR = "ENABLED";
    FD1S3IX count_2638__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i30.GSR = "ENABLED";
    FD1S3IX count_2638__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31902), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638__i31.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27093), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27092), .COUT(n27093), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27091), .COUT(n27092), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27090), .COUT(n27091), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27089), .COUT(n27090), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27088), .COUT(n27089), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26909), .S1(n8065));
    defparam sub_2044_add_2_33.INIT0 = 16'h5555;
    defparam sub_2044_add_2_33.INIT1 = 16'h0000;
    defparam sub_2044_add_2_33.INJECT1_0 = "NO";
    defparam sub_2044_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27087), .COUT(n27088), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27288), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_33.INIT1 = 16'h0000;
    defparam count_2638_add_4_33.INJECT1_0 = "NO";
    defparam count_2638_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27287), .COUT(n27288), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_31.INJECT1_0 = "NO";
    defparam count_2638_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27286), .COUT(n27287), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_29.INJECT1_0 = "NO";
    defparam count_2638_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26908), .COUT(n26909));
    defparam sub_2044_add_2_31.INIT0 = 16'h5999;
    defparam sub_2044_add_2_31.INIT1 = 16'h5999;
    defparam sub_2044_add_2_31.INJECT1_0 = "NO";
    defparam sub_2044_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26907), .COUT(n26908));
    defparam sub_2044_add_2_29.INIT0 = 16'h5999;
    defparam sub_2044_add_2_29.INIT1 = 16'h5999;
    defparam sub_2044_add_2_29.INJECT1_0 = "NO";
    defparam sub_2044_add_2_29.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27285), .COUT(n27286), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_27.INJECT1_0 = "NO";
    defparam count_2638_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27086), .COUT(n27087), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27284), .COUT(n27285), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_25.INJECT1_0 = "NO";
    defparam count_2638_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27085), .COUT(n27086), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26906), .COUT(n26907));
    defparam sub_2044_add_2_27.INIT0 = 16'h5999;
    defparam sub_2044_add_2_27.INIT1 = 16'h5999;
    defparam sub_2044_add_2_27.INJECT1_0 = "NO";
    defparam sub_2044_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27084), .COUT(n27085), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27083), .COUT(n27084), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26905), .COUT(n26906));
    defparam sub_2044_add_2_25.INIT0 = 16'h5999;
    defparam sub_2044_add_2_25.INIT1 = 16'h5999;
    defparam sub_2044_add_2_25.INJECT1_0 = "NO";
    defparam sub_2044_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27283), .COUT(n27284), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_23.INJECT1_0 = "NO";
    defparam count_2638_add_4_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27082), .COUT(n27083), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26904), .COUT(n26905));
    defparam sub_2044_add_2_23.INIT0 = 16'h5999;
    defparam sub_2044_add_2_23.INIT1 = 16'h5999;
    defparam sub_2044_add_2_23.INJECT1_0 = "NO";
    defparam sub_2044_add_2_23.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27282), .COUT(n27283), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_21.INJECT1_0 = "NO";
    defparam count_2638_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27281), .COUT(n27282), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_19.INJECT1_0 = "NO";
    defparam count_2638_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26903), .COUT(n26904));
    defparam sub_2044_add_2_21.INIT0 = 16'h5999;
    defparam sub_2044_add_2_21.INIT1 = 16'h5999;
    defparam sub_2044_add_2_21.INJECT1_0 = "NO";
    defparam sub_2044_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27081), .COUT(n27082), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27280), .COUT(n27281), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_17.INJECT1_0 = "NO";
    defparam count_2638_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27080), .COUT(n27081), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27079), .COUT(n27080), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27078), .COUT(n27079), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27078), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27279), .COUT(n27280), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_15.INJECT1_0 = "NO";
    defparam count_2638_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27278), .COUT(n27279), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_13.INJECT1_0 = "NO";
    defparam count_2638_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27277), .COUT(n27278), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_11.INJECT1_0 = "NO";
    defparam count_2638_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27276), .COUT(n27277), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_9.INJECT1_0 = "NO";
    defparam count_2638_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27275), .COUT(n27276), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_7.INJECT1_0 = "NO";
    defparam count_2638_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27274), .COUT(n27275), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_5.INJECT1_0 = "NO";
    defparam count_2638_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27273), .COUT(n27274), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2638_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2638_add_4_3.INJECT1_0 = "NO";
    defparam count_2638_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2638_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27273), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2638_add_4_1.INIT0 = 16'hF000;
    defparam count_2638_add_4_1.INIT1 = 16'h0555;
    defparam count_2638_add_4_1.INJECT1_0 = "NO";
    defparam count_2638_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26902), .COUT(n26903));
    defparam sub_2044_add_2_19.INIT0 = 16'h5999;
    defparam sub_2044_add_2_19.INIT1 = 16'h5999;
    defparam sub_2044_add_2_19.INJECT1_0 = "NO";
    defparam sub_2044_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26901), .COUT(n26902));
    defparam sub_2044_add_2_17.INIT0 = 16'h5999;
    defparam sub_2044_add_2_17.INIT1 = 16'h5999;
    defparam sub_2044_add_2_17.INJECT1_0 = "NO";
    defparam sub_2044_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26900), .COUT(n26901));
    defparam sub_2044_add_2_15.INIT0 = 16'h5999;
    defparam sub_2044_add_2_15.INIT1 = 16'h5999;
    defparam sub_2044_add_2_15.INJECT1_0 = "NO";
    defparam sub_2044_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2044_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26899), .COUT(n26900));
    defparam sub_2044_add_2_13.INIT0 = 16'h5999;
    defparam sub_2044_add_2_13.INIT1 = 16'h5999;
    defparam sub_2044_add_2_13.INJECT1_0 = "NO";
    defparam sub_2044_add_2_13.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (\read_size[2] , debug_c_c, n13708, 
            n31933, databus, n4168, n31991, \register_addr[0] , n13647, 
            \read_size[0] , n31922, Stepper_X_M0_c_0, n14258, n579, 
            prev_step_clk, step_clk, limit_latched, prev_limit_latched, 
            prev_select, n31951, Stepper_X_Step_c, n27768, \register_addr[1] , 
            GND_net, n34, n31915, n608, n610, n1, \control_reg[7] , 
            n13642, n10962, Stepper_X_En_c, Stepper_X_Dir_c, Stepper_X_M2_c_2, 
            Stepper_X_M1_c_1, read_value, VCC_net, Stepper_X_nFault_c, 
            limit_c_0, n24, n31920, n31904, n16744, n7892, n7926) /* synthesis syn_module_defined=1 */ ;
    output \read_size[2] ;
    input debug_c_c;
    input n13708;
    input n31933;
    input [31:0]databus;
    input n4168;
    input n31991;
    input \register_addr[0] ;
    input n13647;
    output \read_size[0] ;
    input n31922;
    output Stepper_X_M0_c_0;
    input n14258;
    input n579;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    output prev_select;
    input n31951;
    output Stepper_X_Step_c;
    output n27768;
    input \register_addr[1] ;
    input GND_net;
    input n34;
    input n31915;
    input n608;
    input n610;
    input n1;
    output \control_reg[7] ;
    input n13642;
    input n10962;
    output Stepper_X_En_c;
    output Stepper_X_Dir_c;
    output Stepper_X_M2_c_2;
    output Stepper_X_M1_c_1;
    output [31:0]read_value;
    input VCC_net;
    input Stepper_X_nFault_c;
    input limit_c_0;
    input n24;
    input n31920;
    input n31904;
    input n16744;
    output n7892;
    output n7926;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]n224;
    wire [31:0]n4169;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n1_c;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n2, n182, int_step, n1_adj_107, n2_adj_108, n49, n62, 
        n58, n50, n41, n60, n54, n42, n52, n38, n56, n46;
    wire [31:0]n6476;
    
    wire n27189, n27188, n27187, n27186, n27185, n27184, n27183, 
        n27182, n27181, n27180, n27179, n27178, n27177, n27176, 
        n27175, n27174, n1_adj_109, n2_adj_110, n1_adj_111, n2_adj_112, 
        n2_adj_114, n30305, n30306, n30307;
    wire [31:0]n99;
    
    wire n30254, n30255, fault_latched, n30295, n30256, n30293, 
        n30294;
    
    FD1P3AX read_size__i2 (.D(n31933), .SP(n13708), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 mux_1607_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4168), 
         .Z(n4169[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i17_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i31 (.D(n4169[31]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4169[30]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4169[29]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4169[28]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4169[27]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4169[26]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4169[25]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4169[24]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4169[23]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    LUT4 i15076_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_c)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15076_2_lut.init = 16'h2222;
    FD1S3IX steps_reg__i22 (.D(n4169[22]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4169[21]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    LUT4 mux_1913_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1913_Mux_4_i2_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i20 (.D(n4169[20]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4169[19]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4169[18]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4169[17]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4169[16]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4169[15]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4169[14]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4169[13]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4169[12]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4169[11]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4169[10]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4169[9]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4169[8]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4169[7]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4169[6]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4169[5]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4169[4]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4169[3]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4169[2]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4169[1]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1607_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4168), 
         .Z(n4169[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i16_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n13647), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4169[0]), .CK(debug_c_c), .CD(n31991), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n31922), .SP(n13708), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 mux_1607_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4168), 
         .Z(n4169[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i15_3_lut.init = 16'hcaca;
    FD1P3AX control_reg_i1 (.D(n579), .SP(n14258), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13647), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31951), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 mux_1607_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4168), 
         .Z(n4169[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4168), 
         .Z(n4169[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4168), 
         .Z(n4169[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4168), 
         .Z(n4169[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4168), 
         .Z(n4169[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i29_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1607_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4168), 
         .Z(n4169[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4168), 
         .Z(n4169[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4168), 
         .Z(n4169[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i27_3_lut.init = 16'hcaca;
    LUT4 i15077_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1_adj_107)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15077_2_lut.init = 16'h2222;
    LUT4 mux_1607_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4168), 
         .Z(n4169[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1913_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2_adj_108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1913_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27768)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[8]), .B(steps_reg[27]), .C(steps_reg[31]), 
         .D(steps_reg[30]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[15]), .B(n52), .C(n38), .D(steps_reg[11]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[20]), .B(steps_reg[18]), .C(steps_reg[24]), 
         .D(steps_reg[4]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[9]), .B(steps_reg[12]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[5]), .B(n56), .C(n46), .D(steps_reg[6]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[7]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[16]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[17]), .B(steps_reg[21]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[19]), .B(steps_reg[3]), .C(steps_reg[22]), 
         .D(steps_reg[13]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[10]), .B(steps_reg[14]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[29]), .B(steps_reg[0]), .C(steps_reg[2]), 
         .D(steps_reg[1]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[28]), .B(steps_reg[23]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1607_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4168), 
         .Z(n4169[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4168), .Z(n4169[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i10_3_lut.init = 16'hcaca;
    PFUMX mux_1913_Mux_3_i3 (.BLUT(n1_adj_107), .ALUT(n2_adj_108), .C0(\register_addr[1] ), 
          .Z(n6476[3]));
    LUT4 mux_1607_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4168), .Z(n4169[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4168), .Z(n4169[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i8_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27189), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27188), .COUT(n27189), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    LUT4 mux_1607_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4168), 
         .Z(n4169[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i25_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27187), .COUT(n27188), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27186), .COUT(n27187), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    LUT4 mux_1607_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4168), .Z(n4169[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i7_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27185), .COUT(n27186), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    LUT4 mux_1607_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4168), .Z(n4169[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i6_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27184), .COUT(n27185), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27183), .COUT(n27184), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    LUT4 mux_1607_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4168), .Z(n4169[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i5_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27182), .COUT(n27183), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27181), .COUT(n27182), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    LUT4 mux_1607_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4168), .Z(n4169[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4168), 
         .Z(n4169[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4168), .Z(n4169[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4168), .Z(n4169[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i2_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27180), .COUT(n27181), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27179), .COUT(n27180), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    LUT4 mux_1607_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4168), 
         .Z(n4169[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i23_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27178), .COUT(n27179), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    PFUMX mux_1913_Mux_4_i3 (.BLUT(n1_c), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n6476[4]));
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27177), .COUT(n27178), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27176), .COUT(n27177), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27175), .COUT(n27176), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 mux_1607_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4168), 
         .Z(n4169[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i22_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27174), .COUT(n27175), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n34), .D1(prev_step_clk), 
          .COUT(n27174), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_1607_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4168), 
         .Z(n4169[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i21_3_lut.init = 16'hcaca;
    PFUMX mux_1913_Mux_5_i3 (.BLUT(n1_adj_109), .ALUT(n2_adj_110), .C0(\register_addr[1] ), 
          .Z(n6476[5]));
    LUT4 mux_1607_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4168), 
         .Z(n4169[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4168), 
         .Z(n4169[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i19_3_lut.init = 16'hcaca;
    PFUMX mux_1913_Mux_6_i3 (.BLUT(n1_adj_111), .ALUT(n2_adj_112), .C0(\register_addr[1] ), 
          .Z(n6476[6]));
    LUT4 mux_1607_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4168), 
         .Z(n4169[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i18_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n31915), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n31915), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n31915), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n31915), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n31915), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n31915), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n31915), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n31915), .PD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n13647), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n13647), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    PFUMX mux_1913_Mux_7_i3 (.BLUT(n1), .ALUT(n2_adj_114), .C0(\register_addr[1] ), 
          .Z(n6476[7]));
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13642), .CD(n10962), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13642), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13642), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n14258), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13642), .PD(n31991), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n14258), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13642), .PD(n31991), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    PFUMX i22897 (.BLUT(n30305), .ALUT(n30306), .C0(\register_addr[1] ), 
          .Z(n30307));
    LUT4 i15075_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_109)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15075_2_lut.init = 16'h2222;
    LUT4 mux_1913_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2_adj_110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1913_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 i15089_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n99[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15089_4_lut.init = 16'hc088;
    LUT4 i14966_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n99[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14966_4_lut.init = 16'hc088;
    LUT4 i14965_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n99[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14965_4_lut.init = 16'hc088;
    LUT4 i14964_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n99[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14964_4_lut.init = 16'hc088;
    LUT4 i14963_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n99[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14963_4_lut.init = 16'hc088;
    LUT4 i14962_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n99[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14962_4_lut.init = 16'hc088;
    LUT4 i14961_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n99[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14961_4_lut.init = 16'hc088;
    LUT4 i14960_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n99[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14960_4_lut.init = 16'hc088;
    LUT4 i14959_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n99[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14959_4_lut.init = 16'hc088;
    LUT4 i14956_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n99[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14956_4_lut.init = 16'hc088;
    LUT4 i14955_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n99[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14955_4_lut.init = 16'hc088;
    LUT4 i14954_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n99[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14954_4_lut.init = 16'hc088;
    LUT4 i14953_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n99[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14953_4_lut.init = 16'hc088;
    LUT4 i14952_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n99[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14952_4_lut.init = 16'hc088;
    LUT4 i15152_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n99[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15152_4_lut.init = 16'hc088;
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[16]), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n99[16])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i15182_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n99[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15182_4_lut.init = 16'hc088;
    LUT4 i15181_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n99[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15181_4_lut.init = 16'hc088;
    LUT4 i15180_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n99[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15180_4_lut.init = 16'hc088;
    LUT4 i15177_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n99[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15177_4_lut.init = 16'hc088;
    LUT4 i15176_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n99[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15176_4_lut.init = 16'hc088;
    LUT4 i15175_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n99[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15175_4_lut.init = 16'hc088;
    LUT4 i15174_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n99[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15174_4_lut.init = 16'hc088;
    LUT4 i15171_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n99[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15171_4_lut.init = 16'hc088;
    LUT4 i15074_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_111)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15074_2_lut.init = 16'h2222;
    LUT4 mux_1913_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1913_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 i22844_3_lut (.A(Stepper_X_M0_c_0), .B(div_factor_reg[0]), .C(\register_addr[1] ), 
         .Z(n30254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22844_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4168), .Z(n4169[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i1_3_lut.init = 16'hcaca;
    LUT4 i22845_3_lut (.A(limit_latched), .B(steps_reg[0]), .C(\register_addr[1] ), 
         .Z(n30255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22845_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i31 (.D(n99[31]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n99[30]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n99[29]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n99[28]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n99[27]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n99[26]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n99[25]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n99[24]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n99[23]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n99[22]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n99[21]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n99[20]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n99[19]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n99[18]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n99[17]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n99[16]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n99[15]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n99[14]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n99[13]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n99[12]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n99[11]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n99[10]), .SP(n13708), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n99[9]), .SP(n13708), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n99[8]), .SP(n13708), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6476[7]), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6476[6]), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6476[5]), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6476[4]), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6476[3]), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30307), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30295), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    FD1P3AX int_step_182 (.D(n31920), .SP(n24), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n30256), .SP(n13708), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i22895_3_lut (.A(Stepper_X_M2_c_2), .B(n34), .C(\register_addr[0] ), 
         .Z(n30305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22895_3_lut.init = 16'hcaca;
    LUT4 i22896_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22896_3_lut.init = 16'hcaca;
    PFUMX i22885 (.BLUT(n30293), .ALUT(n30294), .C0(\register_addr[1] ), 
          .Z(n30295));
    LUT4 i22883_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22883_3_lut.init = 16'hcaca;
    LUT4 i22884_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22884_3_lut.init = 16'hcaca;
    LUT4 mux_1913_Mux_7_i2_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), 
         .C(\register_addr[0] ), .Z(n2_adj_114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1913_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4168), 
         .Z(n4169[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1607_i32_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n13647), .CD(n31991), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=584, LSE_RLINE=597 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    PFUMX i22846 (.BLUT(n30254), .ALUT(n30255), .C0(\register_addr[0] ), 
          .Z(n30256));
    ClockDivider_U8 step_clk_gen (.div_factor_reg({div_factor_reg}), .GND_net(GND_net), 
            .step_clk(step_clk), .debug_c_c(debug_c_c), .n31991(n31991), 
            .n31904(n31904), .n16744(n16744), .n7892(n7892), .n7926(n7926)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (div_factor_reg, GND_net, step_clk, debug_c_c, 
            n31991, n31904, n16744, n7892, n7926) /* synthesis syn_module_defined=1 */ ;
    input [31:0]div_factor_reg;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31991;
    input n31904;
    input n16744;
    output n7892;
    output n7926;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26969, n26970, n26968, n26967, n26966, n26965, n26964, 
        n26963, n26962, n26961, n26960, n26959, n26958, n7857;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27363, n27362, n27361, n27360, n27359, n27358, n27357, 
        n27356, n27355, n27354, n27353, n27352, n27351, n27350, 
        n27349, n27348;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n27125;
    wire [31:0]n40;
    
    wire n27124, n27005, n27004, n27123, n27122, n27003, n27121, 
        n27120, n27119, n27118, n27117, n27116, n27002, n27115, 
        n27001, n27000, n26999, n26998, n26997, n27114, n26996, 
        n26995, n27113, n27112, n27111, n27110, n26994, n26993, 
        n26992, n26991, n26990, n26989, n26988, n26987, n26986, 
        n26985, n26984, n26983, n26982, n26981, n26980, n26979, 
        n26978, n26977, n26976, n26975, n26974, n26973, n26972, 
        n26971;
    
    CCU2D sub_2037_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26969), .COUT(n26970));
    defparam sub_2037_add_2_25.INIT0 = 16'hf555;
    defparam sub_2037_add_2_25.INIT1 = 16'hf555;
    defparam sub_2037_add_2_25.INJECT1_0 = "NO";
    defparam sub_2037_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26968), .COUT(n26969));
    defparam sub_2037_add_2_23.INIT0 = 16'hf555;
    defparam sub_2037_add_2_23.INIT1 = 16'hf555;
    defparam sub_2037_add_2_23.INJECT1_0 = "NO";
    defparam sub_2037_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26967), .COUT(n26968));
    defparam sub_2037_add_2_21.INIT0 = 16'hf555;
    defparam sub_2037_add_2_21.INIT1 = 16'hf555;
    defparam sub_2037_add_2_21.INJECT1_0 = "NO";
    defparam sub_2037_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26966), .COUT(n26967));
    defparam sub_2037_add_2_19.INIT0 = 16'hf555;
    defparam sub_2037_add_2_19.INIT1 = 16'hf555;
    defparam sub_2037_add_2_19.INJECT1_0 = "NO";
    defparam sub_2037_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26965), .COUT(n26966));
    defparam sub_2037_add_2_17.INIT0 = 16'hf555;
    defparam sub_2037_add_2_17.INIT1 = 16'hf555;
    defparam sub_2037_add_2_17.INJECT1_0 = "NO";
    defparam sub_2037_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26964), .COUT(n26965));
    defparam sub_2037_add_2_15.INIT0 = 16'hf555;
    defparam sub_2037_add_2_15.INIT1 = 16'hf555;
    defparam sub_2037_add_2_15.INJECT1_0 = "NO";
    defparam sub_2037_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26963), .COUT(n26964));
    defparam sub_2037_add_2_13.INIT0 = 16'hf555;
    defparam sub_2037_add_2_13.INIT1 = 16'hf555;
    defparam sub_2037_add_2_13.INJECT1_0 = "NO";
    defparam sub_2037_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26962), .COUT(n26963));
    defparam sub_2037_add_2_11.INIT0 = 16'hf555;
    defparam sub_2037_add_2_11.INIT1 = 16'hf555;
    defparam sub_2037_add_2_11.INJECT1_0 = "NO";
    defparam sub_2037_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26961), .COUT(n26962));
    defparam sub_2037_add_2_9.INIT0 = 16'hf555;
    defparam sub_2037_add_2_9.INIT1 = 16'hf555;
    defparam sub_2037_add_2_9.INJECT1_0 = "NO";
    defparam sub_2037_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26960), .COUT(n26961));
    defparam sub_2037_add_2_7.INIT0 = 16'hf555;
    defparam sub_2037_add_2_7.INIT1 = 16'hf555;
    defparam sub_2037_add_2_7.INJECT1_0 = "NO";
    defparam sub_2037_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26959), .COUT(n26960));
    defparam sub_2037_add_2_5.INIT0 = 16'hf555;
    defparam sub_2037_add_2_5.INIT1 = 16'hf555;
    defparam sub_2037_add_2_5.INJECT1_0 = "NO";
    defparam sub_2037_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26958), .COUT(n26959));
    defparam sub_2037_add_2_3.INIT0 = 16'hf555;
    defparam sub_2037_add_2_3.INIT1 = 16'hf555;
    defparam sub_2037_add_2_3.INJECT1_0 = "NO";
    defparam sub_2037_add_2_3.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7857), .CK(debug_c_c), .CD(n31991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2037_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26958));
    defparam sub_2037_add_2_1.INIT0 = 16'h0000;
    defparam sub_2037_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2037_add_2_1.INJECT1_0 = "NO";
    defparam sub_2037_add_2_1.INJECT1_1 = "NO";
    FD1S3IX count_2636__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i0.GSR = "ENABLED";
    CCU2D count_2636_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27363), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_33.INIT1 = 16'h0000;
    defparam count_2636_add_4_33.INJECT1_0 = "NO";
    defparam count_2636_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27362), .COUT(n27363), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_31.INJECT1_0 = "NO";
    defparam count_2636_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27361), .COUT(n27362), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_29.INJECT1_0 = "NO";
    defparam count_2636_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27360), .COUT(n27361), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_27.INJECT1_0 = "NO";
    defparam count_2636_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27359), .COUT(n27360), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_25.INJECT1_0 = "NO";
    defparam count_2636_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27358), .COUT(n27359), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_23.INJECT1_0 = "NO";
    defparam count_2636_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27357), .COUT(n27358), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_21.INJECT1_0 = "NO";
    defparam count_2636_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27356), .COUT(n27357), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_19.INJECT1_0 = "NO";
    defparam count_2636_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27355), .COUT(n27356), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_17.INJECT1_0 = "NO";
    defparam count_2636_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27354), .COUT(n27355), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_15.INJECT1_0 = "NO";
    defparam count_2636_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27353), .COUT(n27354), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_13.INJECT1_0 = "NO";
    defparam count_2636_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27352), .COUT(n27353), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_11.INJECT1_0 = "NO";
    defparam count_2636_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27351), .COUT(n27352), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_9.INJECT1_0 = "NO";
    defparam count_2636_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27350), .COUT(n27351), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_7.INJECT1_0 = "NO";
    defparam count_2636_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27349), .COUT(n27350), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_5.INJECT1_0 = "NO";
    defparam count_2636_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27348), .COUT(n27349), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2636_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2636_add_4_3.INJECT1_0 = "NO";
    defparam count_2636_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2636_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27348), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636_add_4_1.INIT0 = 16'hF000;
    defparam count_2636_add_4_1.INIT1 = 16'h0555;
    defparam count_2636_add_4_1.INJECT1_0 = "NO";
    defparam count_2636_add_4_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31904), .PD(n16744), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27125), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27124), .COUT(n27125), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27005), .S1(n7857));
    defparam sub_2034_add_2_33.INIT0 = 16'h5555;
    defparam sub_2034_add_2_33.INIT1 = 16'h0000;
    defparam sub_2034_add_2_33.INJECT1_0 = "NO";
    defparam sub_2034_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27004), .COUT(n27005));
    defparam sub_2034_add_2_31.INIT0 = 16'h5999;
    defparam sub_2034_add_2_31.INIT1 = 16'h5999;
    defparam sub_2034_add_2_31.INJECT1_0 = "NO";
    defparam sub_2034_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27123), .COUT(n27124), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27122), .COUT(n27123), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27003), .COUT(n27004));
    defparam sub_2034_add_2_29.INIT0 = 16'h5999;
    defparam sub_2034_add_2_29.INIT1 = 16'h5999;
    defparam sub_2034_add_2_29.INJECT1_0 = "NO";
    defparam sub_2034_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27121), .COUT(n27122), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27120), .COUT(n27121), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27119), .COUT(n27120), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27118), .COUT(n27119), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27117), .COUT(n27118), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27116), .COUT(n27117), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    FD1S3IX count_2636__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i1.GSR = "ENABLED";
    CCU2D sub_2034_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27002), .COUT(n27003));
    defparam sub_2034_add_2_27.INIT0 = 16'h5999;
    defparam sub_2034_add_2_27.INIT1 = 16'h5999;
    defparam sub_2034_add_2_27.INJECT1_0 = "NO";
    defparam sub_2034_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27115), .COUT(n27116), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27001), .COUT(n27002));
    defparam sub_2034_add_2_25.INIT0 = 16'h5999;
    defparam sub_2034_add_2_25.INIT1 = 16'h5999;
    defparam sub_2034_add_2_25.INJECT1_0 = "NO";
    defparam sub_2034_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27000), .COUT(n27001));
    defparam sub_2034_add_2_23.INIT0 = 16'h5999;
    defparam sub_2034_add_2_23.INIT1 = 16'h5999;
    defparam sub_2034_add_2_23.INJECT1_0 = "NO";
    defparam sub_2034_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26999), .COUT(n27000));
    defparam sub_2034_add_2_21.INIT0 = 16'h5999;
    defparam sub_2034_add_2_21.INIT1 = 16'h5999;
    defparam sub_2034_add_2_21.INJECT1_0 = "NO";
    defparam sub_2034_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26998), .COUT(n26999));
    defparam sub_2034_add_2_19.INIT0 = 16'h5999;
    defparam sub_2034_add_2_19.INIT1 = 16'h5999;
    defparam sub_2034_add_2_19.INJECT1_0 = "NO";
    defparam sub_2034_add_2_19.INJECT1_1 = "NO";
    FD1S3IX count_2636__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i2.GSR = "ENABLED";
    FD1S3IX count_2636__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i3.GSR = "ENABLED";
    FD1S3IX count_2636__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i4.GSR = "ENABLED";
    FD1S3IX count_2636__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i5.GSR = "ENABLED";
    FD1S3IX count_2636__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i6.GSR = "ENABLED";
    FD1S3IX count_2636__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i7.GSR = "ENABLED";
    FD1S3IX count_2636__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i8.GSR = "ENABLED";
    FD1S3IX count_2636__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i9.GSR = "ENABLED";
    FD1S3IX count_2636__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i10.GSR = "ENABLED";
    FD1S3IX count_2636__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i11.GSR = "ENABLED";
    FD1S3IX count_2636__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i12.GSR = "ENABLED";
    FD1S3IX count_2636__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i13.GSR = "ENABLED";
    FD1S3IX count_2636__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i14.GSR = "ENABLED";
    FD1S3IX count_2636__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i15.GSR = "ENABLED";
    FD1S3IX count_2636__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i16.GSR = "ENABLED";
    FD1S3IX count_2636__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i17.GSR = "ENABLED";
    FD1S3IX count_2636__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i18.GSR = "ENABLED";
    FD1S3IX count_2636__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i19.GSR = "ENABLED";
    FD1S3IX count_2636__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i20.GSR = "ENABLED";
    FD1S3IX count_2636__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i21.GSR = "ENABLED";
    FD1S3IX count_2636__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i22.GSR = "ENABLED";
    FD1S3IX count_2636__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i23.GSR = "ENABLED";
    FD1S3IX count_2636__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i24.GSR = "ENABLED";
    FD1S3IX count_2636__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i25.GSR = "ENABLED";
    FD1S3IX count_2636__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i26.GSR = "ENABLED";
    FD1S3IX count_2636__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i27.GSR = "ENABLED";
    FD1S3IX count_2636__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i28.GSR = "ENABLED";
    FD1S3IX count_2636__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i29.GSR = "ENABLED";
    FD1S3IX count_2636__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i30.GSR = "ENABLED";
    FD1S3IX count_2636__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31904), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2636__i31.GSR = "ENABLED";
    CCU2D sub_2034_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26997), .COUT(n26998));
    defparam sub_2034_add_2_17.INIT0 = 16'h5999;
    defparam sub_2034_add_2_17.INIT1 = 16'h5999;
    defparam sub_2034_add_2_17.INJECT1_0 = "NO";
    defparam sub_2034_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27114), .COUT(n27115), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26996), .COUT(n26997));
    defparam sub_2034_add_2_15.INIT0 = 16'h5999;
    defparam sub_2034_add_2_15.INIT1 = 16'h5999;
    defparam sub_2034_add_2_15.INJECT1_0 = "NO";
    defparam sub_2034_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26995), .COUT(n26996));
    defparam sub_2034_add_2_13.INIT0 = 16'h5999;
    defparam sub_2034_add_2_13.INIT1 = 16'h5999;
    defparam sub_2034_add_2_13.INJECT1_0 = "NO";
    defparam sub_2034_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27113), .COUT(n27114), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27112), .COUT(n27113), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27111), .COUT(n27112), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27110), .COUT(n27111), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31904), .CD(n16744), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27110), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26994), .COUT(n26995));
    defparam sub_2034_add_2_11.INIT0 = 16'h5999;
    defparam sub_2034_add_2_11.INIT1 = 16'h5999;
    defparam sub_2034_add_2_11.INJECT1_0 = "NO";
    defparam sub_2034_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26993), .COUT(n26994));
    defparam sub_2034_add_2_9.INIT0 = 16'h5999;
    defparam sub_2034_add_2_9.INIT1 = 16'h5999;
    defparam sub_2034_add_2_9.INJECT1_0 = "NO";
    defparam sub_2034_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26992), .COUT(n26993));
    defparam sub_2034_add_2_7.INIT0 = 16'h5999;
    defparam sub_2034_add_2_7.INIT1 = 16'h5999;
    defparam sub_2034_add_2_7.INJECT1_0 = "NO";
    defparam sub_2034_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26991), .COUT(n26992));
    defparam sub_2034_add_2_5.INIT0 = 16'h5999;
    defparam sub_2034_add_2_5.INIT1 = 16'h5999;
    defparam sub_2034_add_2_5.INJECT1_0 = "NO";
    defparam sub_2034_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26990), .COUT(n26991));
    defparam sub_2034_add_2_3.INIT0 = 16'h5999;
    defparam sub_2034_add_2_3.INIT1 = 16'h5999;
    defparam sub_2034_add_2_3.INJECT1_0 = "NO";
    defparam sub_2034_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2034_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26990));
    defparam sub_2034_add_2_1.INIT0 = 16'h0000;
    defparam sub_2034_add_2_1.INIT1 = 16'h5999;
    defparam sub_2034_add_2_1.INJECT1_0 = "NO";
    defparam sub_2034_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26989), .S1(n7892));
    defparam sub_2036_add_2_33.INIT0 = 16'h5999;
    defparam sub_2036_add_2_33.INIT1 = 16'h0000;
    defparam sub_2036_add_2_33.INJECT1_0 = "NO";
    defparam sub_2036_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26988), .COUT(n26989));
    defparam sub_2036_add_2_31.INIT0 = 16'h5999;
    defparam sub_2036_add_2_31.INIT1 = 16'h5999;
    defparam sub_2036_add_2_31.INJECT1_0 = "NO";
    defparam sub_2036_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26987), .COUT(n26988));
    defparam sub_2036_add_2_29.INIT0 = 16'h5999;
    defparam sub_2036_add_2_29.INIT1 = 16'h5999;
    defparam sub_2036_add_2_29.INJECT1_0 = "NO";
    defparam sub_2036_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26986), .COUT(n26987));
    defparam sub_2036_add_2_27.INIT0 = 16'h5999;
    defparam sub_2036_add_2_27.INIT1 = 16'h5999;
    defparam sub_2036_add_2_27.INJECT1_0 = "NO";
    defparam sub_2036_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26985), .COUT(n26986));
    defparam sub_2036_add_2_25.INIT0 = 16'h5999;
    defparam sub_2036_add_2_25.INIT1 = 16'h5999;
    defparam sub_2036_add_2_25.INJECT1_0 = "NO";
    defparam sub_2036_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26984), .COUT(n26985));
    defparam sub_2036_add_2_23.INIT0 = 16'h5999;
    defparam sub_2036_add_2_23.INIT1 = 16'h5999;
    defparam sub_2036_add_2_23.INJECT1_0 = "NO";
    defparam sub_2036_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26983), .COUT(n26984));
    defparam sub_2036_add_2_21.INIT0 = 16'h5999;
    defparam sub_2036_add_2_21.INIT1 = 16'h5999;
    defparam sub_2036_add_2_21.INJECT1_0 = "NO";
    defparam sub_2036_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26982), .COUT(n26983));
    defparam sub_2036_add_2_19.INIT0 = 16'h5999;
    defparam sub_2036_add_2_19.INIT1 = 16'h5999;
    defparam sub_2036_add_2_19.INJECT1_0 = "NO";
    defparam sub_2036_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26981), .COUT(n26982));
    defparam sub_2036_add_2_17.INIT0 = 16'h5999;
    defparam sub_2036_add_2_17.INIT1 = 16'h5999;
    defparam sub_2036_add_2_17.INJECT1_0 = "NO";
    defparam sub_2036_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26980), .COUT(n26981));
    defparam sub_2036_add_2_15.INIT0 = 16'h5999;
    defparam sub_2036_add_2_15.INIT1 = 16'h5999;
    defparam sub_2036_add_2_15.INJECT1_0 = "NO";
    defparam sub_2036_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26979), .COUT(n26980));
    defparam sub_2036_add_2_13.INIT0 = 16'h5999;
    defparam sub_2036_add_2_13.INIT1 = 16'h5999;
    defparam sub_2036_add_2_13.INJECT1_0 = "NO";
    defparam sub_2036_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26978), .COUT(n26979));
    defparam sub_2036_add_2_11.INIT0 = 16'h5999;
    defparam sub_2036_add_2_11.INIT1 = 16'h5999;
    defparam sub_2036_add_2_11.INJECT1_0 = "NO";
    defparam sub_2036_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26977), .COUT(n26978));
    defparam sub_2036_add_2_9.INIT0 = 16'h5999;
    defparam sub_2036_add_2_9.INIT1 = 16'h5999;
    defparam sub_2036_add_2_9.INJECT1_0 = "NO";
    defparam sub_2036_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26976), .COUT(n26977));
    defparam sub_2036_add_2_7.INIT0 = 16'h5999;
    defparam sub_2036_add_2_7.INIT1 = 16'h5999;
    defparam sub_2036_add_2_7.INJECT1_0 = "NO";
    defparam sub_2036_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26975), .COUT(n26976));
    defparam sub_2036_add_2_5.INIT0 = 16'h5999;
    defparam sub_2036_add_2_5.INIT1 = 16'h5999;
    defparam sub_2036_add_2_5.INJECT1_0 = "NO";
    defparam sub_2036_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26974), .COUT(n26975));
    defparam sub_2036_add_2_3.INIT0 = 16'h5999;
    defparam sub_2036_add_2_3.INIT1 = 16'h5999;
    defparam sub_2036_add_2_3.INJECT1_0 = "NO";
    defparam sub_2036_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2036_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26974));
    defparam sub_2036_add_2_1.INIT0 = 16'h0000;
    defparam sub_2036_add_2_1.INIT1 = 16'h5999;
    defparam sub_2036_add_2_1.INJECT1_0 = "NO";
    defparam sub_2036_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26973), .S1(n7926));
    defparam sub_2037_add_2_33.INIT0 = 16'hf555;
    defparam sub_2037_add_2_33.INIT1 = 16'h0000;
    defparam sub_2037_add_2_33.INJECT1_0 = "NO";
    defparam sub_2037_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26972), .COUT(n26973));
    defparam sub_2037_add_2_31.INIT0 = 16'hf555;
    defparam sub_2037_add_2_31.INIT1 = 16'hf555;
    defparam sub_2037_add_2_31.INJECT1_0 = "NO";
    defparam sub_2037_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26971), .COUT(n26972));
    defparam sub_2037_add_2_29.INIT0 = 16'hf555;
    defparam sub_2037_add_2_29.INIT1 = 16'hf555;
    defparam sub_2037_add_2_29.INJECT1_0 = "NO";
    defparam sub_2037_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2037_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26970), .COUT(n26971));
    defparam sub_2037_add_2_27.INIT0 = 16'hf555;
    defparam sub_2037_add_2_27.INIT1 = 16'hf555;
    defparam sub_2037_add_2_27.INJECT1_0 = "NO";
    defparam sub_2037_add_2_27.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module EncoderPeripheral
//

module EncoderPeripheral (\read_size[0] , debug_c_c, n14116, n31950, 
            n31986, prev_select, n31990, read_value, \register_addr[0] , 
            \read_size[2] , n5, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
            n13779, n97, \quadB_delayed[2] , \quadA_delayed[1] , GND_net, 
            n31952, n4433, VCC_net, \quadB_delayed[1] , \quadA_delayed[2] ) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n14116;
    input n31950;
    input n31986;
    output prev_select;
    input n31990;
    output [31:0]read_value;
    input \register_addr[0] ;
    output \read_size[2] ;
    input n5;
    input encoder_ra_c;
    input encoder_rb_c;
    input encoder_ri_c;
    input n13779;
    input n97;
    output \quadB_delayed[2] ;
    output \quadA_delayed[1] ;
    input GND_net;
    input n31952;
    output n4433;
    input VCC_net;
    output \quadB_delayed[1] ;
    output \quadA_delayed[2] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n29724, n29735, n29726, n29733, n29734, n29728, n29720, 
        n29730, n29731;
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    wire n29732, n29723, n29737, n29719, n29722, n29725, n29721, 
        n29729, n29718, n29736, n29727;
    wire [31:0]n180;
    
    FD1P3IX read_size__i1 (.D(n31986), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3AX prev_select_126 (.D(n31990), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam prev_select_126.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29724), .SP(n14116), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29735), .SP(n14116), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29726), .SP(n14116), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29733), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29734), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29728), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29720), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29730), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29731), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [7]), 
         .Z(n29724)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_218 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [8]), 
         .Z(n29735)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_218.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_219 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [9]), 
         .Z(n29726)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_219.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_220 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [10]), 
         .Z(n29733)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_220.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_221 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [11]), 
         .Z(n29734)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_221.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_222 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [12]), 
         .Z(n29728)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_222.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_223 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [13]), 
         .Z(n29720)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_223.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_224 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [14]), 
         .Z(n29730)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_224.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_225 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [15]), 
         .Z(n29731)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_225.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_226 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [16]), 
         .Z(n29732)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_226.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_227 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [17]), 
         .Z(n29723)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_227.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_228 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [18]), 
         .Z(n29737)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_228.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_229 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [19]), 
         .Z(n29719)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_229.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_230 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [20]), 
         .Z(n29722)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_230.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_231 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [21]), 
         .Z(n29725)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_231.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_232 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [22]), 
         .Z(n29721)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_232.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_233 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [23]), 
         .Z(n29729)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_233.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_234 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [24]), 
         .Z(n29718)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_234.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_235 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [26]), 
         .Z(n29736)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_235.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_236 (.A(\register_addr[0] ), .B(n31950), .C(\register[1] [0]), 
         .Z(n29727)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_236.init = 16'h2020;
    FD1P3AX read_value__i16 (.D(n29732), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29723), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29737), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29719), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29722), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29725), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29721), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29729), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29718), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29736), .SP(n14116), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n180[31]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n180[30]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n180[29]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n180[28]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n180[27]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n180[25]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n180[6]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n180[5]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n180[4]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n180[3]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n180[2]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n180[1]), .SP(n14116), .CD(n31950), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n5), .SP(n14116), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i14892_2_lut (.A(\register[1] [31]), .B(\register_addr[0] ), .Z(n180[31])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14892_2_lut.init = 16'h8888;
    LUT4 i14893_2_lut (.A(\register[1] [30]), .B(\register_addr[0] ), .Z(n180[30])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14893_2_lut.init = 16'h8888;
    LUT4 i14894_2_lut (.A(\register[1] [29]), .B(\register_addr[0] ), .Z(n180[29])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14894_2_lut.init = 16'h8888;
    LUT4 i14895_2_lut (.A(\register[1] [28]), .B(\register_addr[0] ), .Z(n180[28])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14895_2_lut.init = 16'h8888;
    LUT4 i14896_2_lut (.A(\register[1] [27]), .B(\register_addr[0] ), .Z(n180[27])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14896_2_lut.init = 16'h8888;
    LUT4 i14897_2_lut (.A(\register[1] [25]), .B(\register_addr[0] ), .Z(n180[25])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14897_2_lut.init = 16'h8888;
    LUT4 i14898_2_lut (.A(\register[1] [6]), .B(\register_addr[0] ), .Z(n180[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14898_2_lut.init = 16'h8888;
    LUT4 i14899_2_lut (.A(\register[1] [5]), .B(\register_addr[0] ), .Z(n180[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14899_2_lut.init = 16'h8888;
    LUT4 i14900_2_lut (.A(\register[1] [4]), .B(\register_addr[0] ), .Z(n180[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam i14900_2_lut.init = 16'h8888;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_ra_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n180[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_rb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n180[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_ri_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n180[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i0 (.D(n29727), .SP(n14116), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=686, LSE_RLINE=696 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(73[9] 89[6])
    defparam read_value__i0.GSR = "ENABLED";
    QuadratureDecoder q (.debug_c_c(debug_c_c), .n13779(n13779), .n97(n97), 
            .quadB_delayed({\quadB_delayed[2] , Open_24, Open_25}), .quadA_delayed({Open_26, 
            \quadA_delayed[1] , Open_27}), .GND_net(GND_net), .n31952(n31952), 
            .n4433(n4433), .\register[1] ({\register[1] }), .VCC_net(VCC_net), 
            .encoder_rb_c(encoder_rb_c), .encoder_ra_c(encoder_ra_c), .\quadB_delayed[1] (\quadB_delayed[1] ), 
            .\quadA_delayed[2] (\quadA_delayed[2] )) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(93[20] 97[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder
//

module QuadratureDecoder (debug_c_c, n13779, n97, quadB_delayed, quadA_delayed, 
            GND_net, n31952, n4433, \register[1] , VCC_net, encoder_rb_c, 
            encoder_ra_c, \quadB_delayed[1] , \quadA_delayed[2] ) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n13779;
    input n97;
    output [2:0]quadB_delayed;
    output [2:0]quadA_delayed;
    input GND_net;
    input n31952;
    output n4433;
    output [31:0]\register[1] ;
    input VCC_net;
    input encoder_rb_c;
    input encoder_ra_c;
    output \quadB_delayed[1] ;
    output \quadA_delayed[2] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    
    wire n26828;
    wire [31:0]n4401;
    
    wire n26827, n26826, n26825, n26824, n26823, n26822, n26821, 
        n26820, n26819, n26818, n26817, n26816, n26815, n26814, 
        n26813;
    wire [2:0]quadB_delayed_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    wire [2:0]quadA_delayed_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    FD1P3AX count__i0 (.D(n97), .SP(n13779), .CK(debug_c_c), .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_1701_33 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[30]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[31]), .D1(GND_net), .CIN(n26828), .S0(n4401[30]), 
          .S1(n4401[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_33.INIT0 = 16'h6969;
    defparam add_1701_33.INIT1 = 16'h6969;
    defparam add_1701_33.INJECT1_0 = "NO";
    defparam add_1701_33.INJECT1_1 = "NO";
    FD1P3IX count__i31 (.D(n4401[31]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4401[30]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n4401[29]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n4401[28]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n4401[27]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n4401[26]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n4401[25]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    CCU2D add_1701_31 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[28]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[29]), .D1(GND_net), .CIN(n26827), .COUT(n26828), 
          .S0(n4401[28]), .S1(n4401[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_31.INIT0 = 16'h6969;
    defparam add_1701_31.INIT1 = 16'h6969;
    defparam add_1701_31.INJECT1_0 = "NO";
    defparam add_1701_31.INJECT1_1 = "NO";
    FD1P3IX count__i24 (.D(n4401[24]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n4401[23]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n4401[22]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n4401[21]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n4401[20]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n4401[19]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n4401[18]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n4401[17]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n4401[16]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n4401[15]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n4401[14]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n4401[13]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n4401[12]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n4401[11]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n4401[10]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n4401[9]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n4401[8]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n4401[7]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n4401[6]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n4401[5]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n4401[4]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n4401[3]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n4401[2]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n4401[1]), .SP(n13779), .CD(n31952), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    CCU2D add_1701_29 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[26]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[27]), .D1(GND_net), .CIN(n26826), .COUT(n26827), 
          .S0(n4401[26]), .S1(n4401[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_29.INIT0 = 16'h6969;
    defparam add_1701_29.INIT1 = 16'h6969;
    defparam add_1701_29.INJECT1_0 = "NO";
    defparam add_1701_29.INJECT1_1 = "NO";
    CCU2D add_1701_27 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[24]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[25]), .D1(GND_net), .CIN(n26825), .COUT(n26826), 
          .S0(n4401[24]), .S1(n4401[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_27.INIT0 = 16'h6969;
    defparam add_1701_27.INIT1 = 16'h6969;
    defparam add_1701_27.INJECT1_0 = "NO";
    defparam add_1701_27.INJECT1_1 = "NO";
    CCU2D add_1701_25 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[22]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[23]), .D1(GND_net), .CIN(n26824), .COUT(n26825), 
          .S0(n4401[22]), .S1(n4401[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_25.INIT0 = 16'h6969;
    defparam add_1701_25.INIT1 = 16'h6969;
    defparam add_1701_25.INJECT1_0 = "NO";
    defparam add_1701_25.INJECT1_1 = "NO";
    CCU2D add_1701_23 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[20]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[21]), .D1(GND_net), .CIN(n26823), .COUT(n26824), 
          .S0(n4401[20]), .S1(n4401[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_23.INIT0 = 16'h6969;
    defparam add_1701_23.INIT1 = 16'h6969;
    defparam add_1701_23.INJECT1_0 = "NO";
    defparam add_1701_23.INJECT1_1 = "NO";
    CCU2D add_1701_21 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[18]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[19]), .D1(GND_net), .CIN(n26822), .COUT(n26823), 
          .S0(n4401[18]), .S1(n4401[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_21.INIT0 = 16'h6969;
    defparam add_1701_21.INIT1 = 16'h6969;
    defparam add_1701_21.INJECT1_0 = "NO";
    defparam add_1701_21.INJECT1_1 = "NO";
    CCU2D add_1701_19 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[16]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[17]), .D1(GND_net), .CIN(n26821), .COUT(n26822), 
          .S0(n4401[16]), .S1(n4401[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_19.INIT0 = 16'h6969;
    defparam add_1701_19.INIT1 = 16'h6969;
    defparam add_1701_19.INJECT1_0 = "NO";
    defparam add_1701_19.INJECT1_1 = "NO";
    CCU2D add_1701_17 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[14]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[15]), .D1(GND_net), .CIN(n26820), .COUT(n26821), 
          .S0(n4401[14]), .S1(n4401[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_17.INIT0 = 16'h6969;
    defparam add_1701_17.INIT1 = 16'h6969;
    defparam add_1701_17.INJECT1_0 = "NO";
    defparam add_1701_17.INJECT1_1 = "NO";
    CCU2D add_1701_15 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[12]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[13]), .D1(GND_net), .CIN(n26819), .COUT(n26820), 
          .S0(n4401[12]), .S1(n4401[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_15.INIT0 = 16'h6969;
    defparam add_1701_15.INIT1 = 16'h6969;
    defparam add_1701_15.INJECT1_0 = "NO";
    defparam add_1701_15.INJECT1_1 = "NO";
    CCU2D add_1701_13 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[10]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[11]), .D1(GND_net), .CIN(n26818), .COUT(n26819), 
          .S0(n4401[10]), .S1(n4401[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_13.INIT0 = 16'h6969;
    defparam add_1701_13.INIT1 = 16'h6969;
    defparam add_1701_13.INJECT1_0 = "NO";
    defparam add_1701_13.INJECT1_1 = "NO";
    CCU2D add_1701_11 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[8]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[9]), .D1(GND_net), .CIN(n26817), .COUT(n26818), 
          .S0(n4401[8]), .S1(n4401[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_11.INIT0 = 16'h6969;
    defparam add_1701_11.INIT1 = 16'h6969;
    defparam add_1701_11.INJECT1_0 = "NO";
    defparam add_1701_11.INJECT1_1 = "NO";
    CCU2D add_1701_9 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[6]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[7]), .D1(GND_net), .CIN(n26816), .COUT(n26817), 
          .S0(n4401[6]), .S1(n4401[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_9.INIT0 = 16'h6969;
    defparam add_1701_9.INIT1 = 16'h6969;
    defparam add_1701_9.INJECT1_0 = "NO";
    defparam add_1701_9.INJECT1_1 = "NO";
    CCU2D add_1701_7 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[4]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[5]), .D1(GND_net), .CIN(n26815), .COUT(n26816), 
          .S0(n4401[4]), .S1(n4401[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_7.INIT0 = 16'h6969;
    defparam add_1701_7.INIT1 = 16'h6969;
    defparam add_1701_7.INJECT1_0 = "NO";
    defparam add_1701_7.INJECT1_1 = "NO";
    CCU2D add_1701_5 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[2]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[3]), .D1(GND_net), .CIN(n26814), .COUT(n26815), 
          .S0(n4401[2]), .S1(n4401[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_5.INIT0 = 16'h6969;
    defparam add_1701_5.INIT1 = 16'h6969;
    defparam add_1701_5.INJECT1_0 = "NO";
    defparam add_1701_5.INJECT1_1 = "NO";
    CCU2D add_1701_3 (.A0(quadB_delayed[2]), .B0(quadA_delayed[1]), .C0(count[0]), 
          .D0(GND_net), .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), 
          .C1(count[1]), .D1(GND_net), .CIN(n26813), .COUT(n26814), 
          .S0(n4433), .S1(n4401[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_3.INIT0 = 16'h9696;
    defparam add_1701_3.INIT1 = 16'h6969;
    defparam add_1701_3.INJECT1_0 = "NO";
    defparam add_1701_3.INJECT1_1 = "NO";
    CCU2D add_1701_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quadB_delayed[2]), .B1(quadA_delayed[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26813));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1701_1.INIT0 = 16'hF000;
    defparam add_1701_1.INIT1 = 16'h6666;
    defparam add_1701_1.INJECT1_0 = "NO";
    defparam add_1701_1.INJECT1_1 = "NO";
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_rb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed_c[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_ra_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed_c[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(n31952), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed_c[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed_c[0]), .CK(debug_c_c), .Q(quadA_delayed[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(quadA_delayed[1]), .CK(debug_c_c), .Q(\quadA_delayed[2] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=93, LSE_RLINE=97 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (databus, register_addr, n32090, 
            n30166, debug_c_c, \select[7] , n31975, n32001, prev_select, 
            n31923, \select[4] , \select[3] , \select[2] , \select[1] , 
            databus_out, n13608, n32075, rw, n31926, n1486, debug_c_7, 
            n31928, n31911, n224, n3899, prev_select_adj_1, n31991, 
            n13876, \sendcount[1] , n32052, n8, n31944, n32032, 
            n32089, n29768, n32011, n29174, n29175, n31996, n31965, 
            \read_value[1] , n4, n13700, n31972, n29770, n32056, 
            n11158, prev_select_adj_2, n31986, \read_value[28] , n33683, 
            n3, n27768, \control_reg[7] , n32088, n34, n31933, n29916, 
            n13647, n32005, \register[2][3] , n5980, n27787, \control_reg[7]_adj_3 , 
            n32, prev_select_adj_4, n27886, n33682, n13323, n31938, 
            \read_value[27] , n3_adj_5, n29798, n31937, n33680, n15, 
            n31940, n250_adj_6, n32034, n31982, n31955, n4071, n13708, 
            n32003, n94, n32006, \register[2][4] , n29197, \register[2][5] , 
            n29211, \register[2][6] , n29213, \register[2][7] , n29207, 
            \register[2][8] , n29199, \register[2][9] , n29215, \register[2][10] , 
            n29189, n31915, n31990, \register[2][11] , n29190, \register[2][12] , 
            n29201, \register[2][13] , n29209, \register[2][14] , n29203, 
            n14372, n9362, n12930, \register[2][15] , n29191, \register[2][16] , 
            n29193, n22, n12, n8_adj_7, \register[2][17] , n29205, 
            \reg_size[2] , n32068, n32004, n5811, n27946, n31951, 
            n52, \register[2][18] , n29194, n1480, n31977, \register[2][19] , 
            n29196, \register[2][20] , n29198, \register[2][21] , n29200, 
            n1483, \register[2][22] , n29202, \register[2][23] , n29204, 
            n32030, \register[2][24] , n29206, \register[2][25] , n29208, 
            \register[2][26] , n29210, \register[2][27] , n29214, n4_adj_8, 
            \register[2][28] , n29216, \register[2][29] , n29195, \register[2][30] , 
            n29192, \register[2][31] , n29212, n31987, n31953, n14094, 
            n31970, n31910, n13710, \read_value[26] , n3_adj_9, \read_value[25] , 
            n3_adj_10, \read_value[24] , n3_adj_11, \steps_reg[5] , 
            n14, \steps_reg[6] , n13, \steps_reg[3] , n12_adj_12, 
            \read_value[23] , n3_adj_13, \read_value[22] , n3_adj_14, 
            \control_reg[7]_adj_15 , n8494, \read_value[21] , n3_adj_16, 
            \read_value[20] , n3_adj_17, \read_value[19] , n3_adj_18, 
            \read_value[18] , n3_adj_19, n13642, \control_reg[7]_adj_20 , 
            n8476, \read_value[17] , n3_adj_21, \read_value[16] , n3_adj_22, 
            \read_value[15] , n3_adj_23, \read_value[14] , n3_adj_24, 
            n13667, \read_value[13] , n3_adj_25, n3984, \read_value[12] , 
            n3_adj_26, \read_value[11] , n3_adj_27, n13693, n9139, 
            n1, n31942, \read_value[10] , n3_adj_28, \read_value[9] , 
            n3_adj_29, \read_value[8] , n3_adj_30, debug_c_2, debug_c_3, 
            n27766, n32_adj_31, debug_c_4, debug_c_5, n31921, n14661, 
            n31922, n96, \read_value[31] , n3_adj_32, \read_value[29] , 
            n3_adj_33, n8485, \read_value[30] , n3_adj_34, prev_select_adj_35, 
            n5, n27769, n32_adj_36, \reset_count[14] , \reset_count[13] , 
            \reset_count[12] , n29900, n10889, GND_net, uart_rx_c) /* synthesis syn_module_defined=1 */ ;
    input [31:0]databus;
    output [7:0]register_addr;
    output n32090;
    output n30166;
    input debug_c_c;
    output \select[7] ;
    input n31975;
    output n32001;
    input prev_select;
    output n31923;
    output \select[4] ;
    output \select[3] ;
    output \select[2] ;
    output \select[1] ;
    output [31:0]databus_out;
    input n13608;
    input n32075;
    output rw;
    output n31926;
    output n1486;
    output debug_c_7;
    input n31928;
    input n31911;
    input [31:0]n224;
    output [31:0]n3899;
    input prev_select_adj_1;
    input n31991;
    output n13876;
    output \sendcount[1] ;
    output n32052;
    output n8;
    output n31944;
    output n32032;
    output n32089;
    output n29768;
    output n32011;
    output n29174;
    output n29175;
    output n31996;
    input n31965;
    input \read_value[1] ;
    output n4;
    output n13700;
    input n31972;
    output n29770;
    output n32056;
    output n11158;
    input prev_select_adj_2;
    output n31986;
    input \read_value[28] ;
    output n33683;
    output n3;
    input n27768;
    input \control_reg[7] ;
    input n32088;
    output n34;
    output n31933;
    output n29916;
    output n13647;
    output n32005;
    input \register[2][3] ;
    output n5980;
    input n27787;
    input \control_reg[7]_adj_3 ;
    output n32;
    input prev_select_adj_4;
    input n27886;
    input n33682;
    input n13323;
    output n31938;
    input \read_value[27] ;
    output n3_adj_5;
    output n29798;
    output n31937;
    output n33680;
    output n15;
    output n31940;
    output n250_adj_6;
    output n32034;
    output n31982;
    input n31955;
    output n4071;
    output n13708;
    output n32003;
    output n94;
    input n32006;
    input \register[2][4] ;
    output n29197;
    input \register[2][5] ;
    output n29211;
    input \register[2][6] ;
    output n29213;
    input \register[2][7] ;
    output n29207;
    input \register[2][8] ;
    output n29199;
    input \register[2][9] ;
    output n29215;
    input \register[2][10] ;
    output n29189;
    output n31915;
    output n31990;
    input \register[2][11] ;
    output n29190;
    input \register[2][12] ;
    output n29201;
    input \register[2][13] ;
    output n29209;
    input \register[2][14] ;
    output n29203;
    input n14372;
    output n9362;
    input n12930;
    input \register[2][15] ;
    output n29191;
    input \register[2][16] ;
    output n29193;
    input n22;
    input n12;
    input n8_adj_7;
    input \register[2][17] ;
    output n29205;
    input \reg_size[2] ;
    input n32068;
    output n32004;
    output n5811;
    output n27946;
    output n31951;
    output n52;
    input \register[2][18] ;
    output n29194;
    output n1480;
    output n31977;
    input \register[2][19] ;
    output n29196;
    input \register[2][20] ;
    output n29198;
    input \register[2][21] ;
    output n29200;
    output n1483;
    input \register[2][22] ;
    output n29202;
    input \register[2][23] ;
    output n29204;
    output n32030;
    input \register[2][24] ;
    output n29206;
    input \register[2][25] ;
    output n29208;
    input \register[2][26] ;
    output n29210;
    input \register[2][27] ;
    output n29214;
    output n4_adj_8;
    input \register[2][28] ;
    output n29216;
    input \register[2][29] ;
    output n29195;
    input \register[2][30] ;
    output n29192;
    input \register[2][31] ;
    output n29212;
    input n31987;
    output n31953;
    output n14094;
    input n31970;
    output n31910;
    output n13710;
    input \read_value[26] ;
    output n3_adj_9;
    input \read_value[25] ;
    output n3_adj_10;
    input \read_value[24] ;
    output n3_adj_11;
    input \steps_reg[5] ;
    output n14;
    input \steps_reg[6] ;
    output n13;
    input \steps_reg[3] ;
    output n12_adj_12;
    input \read_value[23] ;
    output n3_adj_13;
    input \read_value[22] ;
    output n3_adj_14;
    input \control_reg[7]_adj_15 ;
    output n8494;
    input \read_value[21] ;
    output n3_adj_16;
    input \read_value[20] ;
    output n3_adj_17;
    input \read_value[19] ;
    output n3_adj_18;
    input \read_value[18] ;
    output n3_adj_19;
    output n13642;
    input \control_reg[7]_adj_20 ;
    output n8476;
    input \read_value[17] ;
    output n3_adj_21;
    input \read_value[16] ;
    output n3_adj_22;
    input \read_value[15] ;
    output n3_adj_23;
    input \read_value[14] ;
    output n3_adj_24;
    output n13667;
    input \read_value[13] ;
    output n3_adj_25;
    output n3984;
    input \read_value[12] ;
    output n3_adj_26;
    input \read_value[11] ;
    output n3_adj_27;
    output n13693;
    output n9139;
    output n1;
    output n31942;
    input \read_value[10] ;
    output n3_adj_28;
    input \read_value[9] ;
    output n3_adj_29;
    input \read_value[8] ;
    output n3_adj_30;
    output debug_c_2;
    output debug_c_3;
    input n27766;
    output n32_adj_31;
    output debug_c_4;
    output debug_c_5;
    output n31921;
    output n14661;
    output n31922;
    output n96;
    input \read_value[31] ;
    output n3_adj_32;
    input \read_value[29] ;
    output n3_adj_33;
    output n8485;
    input \read_value[30] ;
    output n3_adj_34;
    input prev_select_adj_35;
    output n5;
    input n27769;
    output n32_adj_36;
    input \reset_count[14] ;
    input \reset_count[13] ;
    input \reset_count[12] ;
    input n29900;
    output n10889;
    input GND_net;
    input uart_rx_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(461[15:21])
    wire n33682 /* synthesis nomerge= */ ;
    
    wire n5_c;
    wire [31:0]n1468;
    
    wire n29688, n27931;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n29972, n5_adj_1, n29691, n27929, n5_adj_2, n29685, n27933, 
        n5_adj_3, n29689, n27927, n5_adj_4, n29681, n27937;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n31971;
    wire [4:0]n18;
    
    wire n33689, n15373, n15377, n31899, n31900, n16362, n2800;
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    wire [7:0]n5802;
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n32099, n32475, n15369;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n31960;
    wire [7:0]n2210;
    
    wire n5_adj_5, n29694, n27885, n15389, n31117, n29971, n2798;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n167, n5_adj_6, n29690, n27928;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n14791, n28838, n13536, n32041, n31229, n31230, n2738, 
        n32042, n30186, n21696, n31984, n5_adj_7, n29693, n27889, 
        n32043, n29185, escape, n32044, n31962, n32045, n32018, 
        n7, n32046, n32021, n32047, n30007, n32048, n6, n32008, 
        n29889, n32094, n31673, n31674, n32098, n32097, n32101, 
        n32100, n32104, n32103, n31675, n5_adj_9, n29692, n27930, 
        n32033, n32078, n32107, n32106, n32110, n32109, n32113, 
        n32112, n32116, n32115, n32119, n32118, n32122, n32121, 
        n31936, n32012, n13148, n6_adj_10, n10796;
    wire [4:0]n19;
    
    wire n5_adj_11, n29695, n27906, n5_adj_12, n29696, n27851, n5_adj_13, 
        n29683, n27870, n32474, n32017, n32472, n32473, n5_adj_14, 
        n29697, n27863, n4_adj_16, n32057, n9_adj_17, n31983, n5_adj_18, 
        n29679, n27862, n29984, n32059, n5_adj_19, n29698, n27852, 
        n32020, n5_adj_20, n29699, n27848, n5_adj_21, n29700, n27897, 
        n32061, n5_adj_22, n29701, n27861, n31115, n5_adj_23, n29702, 
        n27847, n5_adj_24, n29703, n27860, n5_adj_25, n29704, n27849, 
        n5_adj_26, n29705, n27845, n29983, n5_adj_27, n29706, n27836, 
        n5_adj_28, n29707, n27856, n2219, n5_adj_29, n29708, n27855, 
        n13177, send, n5_adj_32, n29709, n27822, n5_adj_33, n29682, 
        n27824, n31111, n7_adj_34, n31118, n30136, n5_adj_36, n29680, 
        n27842, n29904, n5_adj_38, n29710, n27838, n11_adj_39, n11_adj_40, 
        n11_adj_41, n11_adj_42, n11_adj_43, n11_adj_44, n11_adj_45, 
        n11_adj_46, n4_adj_47, n32105;
    wire [7:0]n9241;
    
    wire n4_adj_48, n32108, n4_adj_49, n32111, n4_adj_50, n32117;
    wire [3:0]n1864;
    
    wire n1921, n12_c, n14_c, n28826, n16363, n15376, n15366, 
        n15372, n16361, n29883, n29684, n4_adj_51, n32123, n4_adj_52, 
        n32120, n27964, n28822, n32102, n31116, n4_adj_53, n32114, 
        n13275, n29673, n29981, n29980, n28836, n28858, n28814, 
        n28844, n28842, n11_adj_54, n28834, n29686, n8_adj_55, n29014, 
        n11_adj_56, n28900, n15_adj_57, n29663, n29835, n11_adj_58, 
        n28840, n1_c, n6_adj_59, n11_adj_60, n11_adj_61, n11_adj_62, 
        n11_adj_63, n11_adj_64, n28076, n29922, n28884, n28850, 
        n28824, n29605, n28988, n28916, n30106, n1573, n28818, 
        n2, n29600, n15368, n1869, n5_adj_67, n27934, n15388, 
        busy, n1579, n1580, n5_adj_68, n27872, n5_adj_69, n29687, 
        n27926, n6_adj_70;
    wire [7:0]register_addr_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:26])
    
    wire n11026, n12151, n38, n28948, n31218, n11000, n12261, 
        n12818, n31966, n12149;
    wire [3:0]n9543;
    
    wire n16499, n4_adj_91, n16497, n32095, n10, n29997, n8_adj_98, 
        n8_adj_100, n30102, n29715;
    
    LUT4 i2_4_lut (.A(databus[3]), .B(n5_c), .C(n1468[13]), .D(n29688), 
         .Z(n27931)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 select_2107_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1468[4]), 
         .C(rx_data[3]), .D(n29972), .Z(n5_c)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i22758_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[4]), 
         .C(register_addr[3]), .D(n32090), .Z(n30166)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22758_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_26 (.A(databus[4]), .B(n5_adj_1), .C(n1468[13]), 
         .D(n29691), .Z(n27929)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_26.init = 16'hffec;
    LUT4 select_2107_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1468[4]), 
         .C(rx_data[4]), .D(n29972), .Z(n5_adj_1)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_27 (.A(databus[5]), .B(n5_adj_2), .C(n1468[13]), 
         .D(n29685), .Z(n27933)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_27.init = 16'hffec;
    LUT4 select_2107_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1468[4]), 
         .C(rx_data[5]), .D(n29972), .Z(n5_adj_2)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_28 (.A(databus[6]), .B(n5_adj_3), .C(n1468[13]), 
         .D(n29689), .Z(n27927)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_28.init = 16'hffec;
    LUT4 select_2107_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1468[4]), 
         .C(rx_data[6]), .D(n29972), .Z(n5_adj_3)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_29 (.A(databus[7]), .B(n5_adj_4), .C(n1468[13]), 
         .D(n29681), .Z(n27937)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_29.init = 16'hffec;
    LUT4 select_2107_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1468[4]), 
         .C(rx_data[7]), .D(n29972), .Z(n5_adj_4)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_23_i5_4_lut.init = 16'h88c0;
    FD1P3AX sendcount__i0 (.D(n18[0]), .SP(n31971), .CK(debug_c_c), .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    FD1S3IX select__i7 (.D(n15373), .CK(debug_c_c), .CD(n33689), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_306_4_lut (.A(register_addr[1]), .B(n31975), .C(n32001), 
         .D(prev_select), .Z(n31923)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_306_4_lut.init = 16'h00e0;
    FD1S3IX select__i4 (.D(n15377), .CK(debug_c_c), .CD(n33689), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1S3IX select__i3 (.D(n31899), .CK(debug_c_c), .CD(n33689), .Q(\select[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i3.GSR = "ENABLED";
    FD1S3IX select__i2 (.D(n31900), .CK(debug_c_c), .CD(n33689), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1S3IX select__i1 (.D(n16362), .CK(debug_c_c), .CD(n33689), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i4 (.D(n5802[4]), .SP(n13608), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n5802[2]), .SP(n13608), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n5802[1]), .SP(n13608), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    FD1S3IX bufcount__i3 (.D(n32099), .CK(debug_c_c), .CD(n33689), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n32475), .CK(debug_c_c), .CD(n33689), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n15369), .CK(debug_c_c), .CD(n33689), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2210[4]), .SP(n31960), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_30 (.A(databus[8]), .B(n5_adj_5), .C(n1468[13]), 
         .D(n29694), .Z(n27885)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_30.init = 16'hffec;
    FD1P3AX tx_data_i0_i3 (.D(n2210[3]), .SP(n31960), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n2210[0]), .SP(n31960), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n15389), .CK(debug_c_c), .CD(n33689), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n31117), .SP(n13608), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2800), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2210[1]), .SP(n31960), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_309_4_lut (.A(register_addr[1]), .B(n31975), .C(n32075), 
         .D(rw), .Z(n31926)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_309_4_lut.init = 16'h0010;
    LUT4 select_2107_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1468[4]), 
         .C(rx_data[0]), .D(n29971), .Z(n5_adj_5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_24_i5_4_lut.init = 16'h88c0;
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\select[4] ), .B(register_addr[5]), .Z(n167)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_31 (.A(databus[9]), .B(n5_adj_6), .C(n1468[13]), 
         .D(n29690), .Z(n27928)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_31.init = 16'hffec;
    FD1P3IX buffer_0___i1 (.D(n28838), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    FD1S3JX state_FSM_i1 (.D(n13536), .CK(debug_c_c), .PD(n33689), .Q(n1468[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_424 (.A(n1486), .B(sendcount[4]), .Z(n32041)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_424.init = 16'h2222;
    LUT4 motor_pwm_r_c_bdd_2_lut_23401_3_lut (.A(n1486), .B(sendcount[4]), 
         .C(n31229), .Z(n31230)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam motor_pwm_r_c_bdd_2_lut_23401_3_lut.init = 16'h2020;
    LUT4 select_2107_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1468[4]), 
         .C(rx_data[1]), .D(n29971), .Z(n5_adj_6)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 mux_522_i5_3_lut (.A(n2738), .B(esc_data[4]), .C(n1468[18]), 
         .Z(n2210[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i5_3_lut.init = 16'hcaca;
    LUT4 i22668_2_lut_rep_425 (.A(rx_data[6]), .B(rx_data[7]), .Z(n32042)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22668_2_lut_rep_425.init = 16'heeee;
    LUT4 i22830_3_lut_rep_367_4_lut (.A(rx_data[6]), .B(rx_data[7]), .C(n30186), 
         .D(n21696), .Z(n31984)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22830_3_lut_rep_367_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_32 (.A(databus[10]), .B(n5_adj_7), .C(n1468[13]), 
         .D(n29693), .Z(n27889)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_32.init = 16'hffec;
    LUT4 i1_2_lut_rep_426 (.A(rx_data[5]), .B(rx_data[0]), .Z(n32043)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i1_2_lut_rep_426.init = 16'hbbbb;
    LUT4 i2_3_lut_4_lut (.A(rx_data[5]), .B(rx_data[0]), .C(rx_data[2]), 
         .D(n32042), .Z(n29185)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i2_3_lut_4_lut.init = 16'hfffb;
    LUT4 i923_2_lut_rep_427 (.A(escape), .B(debug_c_7), .Z(n32044)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i923_2_lut_rep_427.init = 16'hbbbb;
    LUT4 i2_3_lut_rep_345_4_lut (.A(escape), .B(debug_c_7), .C(n31984), 
         .D(n1468[4]), .Z(n31962)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_345_4_lut.init = 16'hfffb;
    LUT4 mux_1537_i15_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[14]), 
         .D(n224[14]), .Z(n3899[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_rep_428 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n32045)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_rep_428.init = 16'hecec;
    LUT4 i2_2_lut_rep_401_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1468[4]), .Z(n32018)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_401_4_lut.init = 16'hecff;
    LUT4 i1_2_lut_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1468[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hec00;
    LUT4 i3262_2_lut_rep_429 (.A(bufcount[1]), .B(bufcount[2]), .Z(n32046)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3262_2_lut_rep_429.init = 16'heeee;
    LUT4 i2897_2_lut_rep_404_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n32021)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2897_2_lut_rep_404_3_lut.init = 16'hfefe;
    LUT4 i4_2_lut_rep_430 (.A(n1486), .B(n1468[15]), .Z(n32047)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_430.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(n1486), .B(n1468[15]), .C(n1468[12]), .Z(n30007)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_431 (.A(n1468[7]), .B(n1468[13]), .C(n1468[5]), 
         .Z(n32048)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_431.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_33 (.A(n1468[7]), .B(n1468[13]), .C(n1468[5]), 
         .D(n1468[6]), .Z(n6)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_33.init = 16'hfffe;
    LUT4 select_2107_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1468[4]), 
         .C(rx_data[2]), .D(n29971), .Z(n5_adj_7)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i2_3_lut_4_lut_adj_34 (.A(n32090), .B(n32008), .C(prev_select_adj_1), 
         .D(n31991), .Z(n13876)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_34.init = 16'h0004;
    LUT4 i1_2_lut_adj_35 (.A(\select[4] ), .B(register_addr[4]), .Z(n29889)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_35.init = 16'h2222;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32094)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 sendcount_1__bdd_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(sendcount[3]), 
         .D(sendcount[2]), .Z(n31673)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_1__bdd_4_lut.init = 16'h6aaa;
    LUT4 sendcount_4__bdd_3_lut (.A(sendcount[4]), .B(n31673), .C(\sendcount[1] ), 
         .Z(n31674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut.init = 16'hcaca;
    LUT4 i20111_2_lut_rep_435 (.A(register_addr[4]), .B(register_addr[0]), 
         .Z(n32052)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20111_2_lut_rep_435.init = 16'heeee;
    LUT4 i3_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[0]), .C(\select[1] ), 
         .D(rw), .Z(n8)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0010;
    LUT4 i8740_then_4_lut (.A(bufcount[3]), .B(n1468[0]), .C(n1468[3]), 
         .D(n1468[4]), .Z(n32098)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8740_then_4_lut.init = 16'haaa2;
    LUT4 i8740_else_4_lut (.A(bufcount[3]), .B(n1468[0]), .C(n1468[3]), 
         .D(n1468[4]), .Z(n32097)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8740_else_4_lut.init = 16'h0002;
    LUT4 i23356_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n32101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23356_then_3_lut.init = 16'hcaca;
    LUT4 i23356_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n32100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23356_else_3_lut.init = 16'hcaca;
    LUT4 i22864_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n32104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22864_then_3_lut.init = 16'hcaca;
    LUT4 i22864_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n32103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22864_else_3_lut.init = 16'hcaca;
    LUT4 rx_data_3__bdd_4_lut_23802 (.A(rx_data[3]), .B(rx_data[2]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n31675)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_3__bdd_4_lut_23802.init = 16'h6001;
    LUT4 i2_4_lut_adj_36 (.A(databus[11]), .B(n5_adj_9), .C(n1468[13]), 
         .D(n29692), .Z(n27930)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_36.init = 16'hffec;
    LUT4 i1_2_lut_rep_327_3_lut_4_lut (.A(n32090), .B(n32033), .C(rw), 
         .D(n32078), .Z(n31944)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_327_3_lut_4_lut.init = 16'h1000;
    LUT4 i22867_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n32107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22867_then_3_lut.init = 16'hcaca;
    LUT4 i22867_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n32106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22867_else_3_lut.init = 16'hcaca;
    LUT4 i22870_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n32110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22870_then_3_lut.init = 16'hcaca;
    LUT4 i22870_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n32109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22870_else_3_lut.init = 16'hcaca;
    LUT4 i22873_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n32113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22873_then_3_lut.init = 16'hcaca;
    LUT4 i22873_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n32112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22873_else_3_lut.init = 16'hcaca;
    LUT4 mux_1537_i2_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[1]), 
         .D(n224[1]), .Z(n3899[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_37 (.A(register_addr[1]), .B(n32032), .C(n32089), 
         .D(register_addr[4]), .Z(n29768)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_37.init = 16'h0200;
    LUT4 i22876_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n32116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22876_then_3_lut.init = 16'hcaca;
    LUT4 mux_1537_i9_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[8]), 
         .D(n224[8]), .Z(n3899[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i22876_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n32115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22876_else_3_lut.init = 16'hcaca;
    LUT4 i22879_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n32119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22879_then_3_lut.init = 16'hcaca;
    LUT4 i22879_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n32118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22879_else_3_lut.init = 16'hcaca;
    LUT4 i22882_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n32122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22882_then_3_lut.init = 16'hcaca;
    LUT4 i22882_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n32121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22882_else_3_lut.init = 16'hcaca;
    FD1P3IX sendcount__i4 (.D(n31674), .SP(n31971), .CD(n31936), .CK(debug_c_c), 
            .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 select_2107_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1468[4]), 
         .C(rx_data[3]), .D(n29971), .Z(n5_adj_9)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_394_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .Z(n32011)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_394_3_lut.init = 16'hfefe;
    LUT4 i23057_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .D(n32012), .Z(n29174)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i23057_3_lut_4_lut.init = 16'h0010;
    LUT4 i23054_2_lut_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n32012), .D(register_addr[1]), .Z(n29175)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i23054_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i9381_4_lut (.A(escape), .B(n13148), .C(n6_adj_10), .D(n1468[3]), 
         .Z(n10796)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i9381_4_lut.init = 16'h1aaa;
    LUT4 i2_2_lut (.A(debug_c_7), .B(n31996), .Z(n6_adj_10)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    FD1P3IX sendcount__i3 (.D(n19[3]), .SP(n31971), .CD(n31936), .CK(debug_c_c), 
            .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3IX sendcount__i2 (.D(n19[2]), .SP(n31971), .CD(n31936), .CK(debug_c_c), 
            .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n19[1]), .SP(n31971), .CD(n31936), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 Select_4253_i4_2_lut_4_lut (.A(\select[4] ), .B(rw), .C(n31965), 
         .D(\read_value[1] ), .Z(n4)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam Select_4253_i4_2_lut_4_lut.init = 16'h0800;
    LUT4 i2_4_lut_adj_38 (.A(databus[12]), .B(n5_adj_11), .C(n1468[13]), 
         .D(n29695), .Z(n27906)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_38.init = 16'hffec;
    LUT4 i2_4_lut_adj_39 (.A(n29185), .B(rx_data[4]), .C(rx_data[1]), 
         .D(rx_data[3]), .Z(n13148)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i2_4_lut_adj_39.init = 16'hbfff;
    LUT4 mux_1537_i8_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[7]), 
         .D(n224[7]), .Z(n3899[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1537_i7_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[6]), 
         .D(n224[6]), .Z(n3899[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 select_2107_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1468[4]), 
         .C(rx_data[4]), .D(n29971), .Z(n5_adj_11)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_40 (.A(databus[13]), .B(n5_adj_12), .C(n1468[13]), 
         .D(n29696), .Z(n27851)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_40.init = 16'hffec;
    LUT4 select_2107_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1468[4]), 
         .C(rx_data[5]), .D(n29971), .Z(n5_adj_12)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_29_i5_4_lut.init = 16'h88c0;
    FD1P3AX rw_498 (.D(n1468[10]), .SP(n2798), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_41 (.A(databus[14]), .B(n5_adj_13), .C(n1468[13]), 
         .D(n29683), .Z(n27870)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_41.init = 16'hffec;
    LUT4 mux_1537_i6_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[5]), 
         .D(n224[5]), .Z(n3899[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_42 (.A(register_addr[4]), .B(n13700), .C(n31972), 
         .D(register_addr[1]), .Z(n29770)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A (B+!(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_42.init = 16'h3b00;
    LUT4 i1_2_lut_rep_439 (.A(register_addr[1]), .B(register_addr[0]), .Z(n32056)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_439.init = 16'heeee;
    LUT4 n31984_bdd_4_lut (.A(bufcount[1]), .B(n1468[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n32474)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n31984_bdd_4_lut.init = 16'h0080;
    FD1S3AX escape_501 (.D(n10796), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 select_2107_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1468[4]), 
         .C(rx_data[6]), .D(n29971), .Z(n5_adj_13)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i260_2_lut_rep_400_3_lut (.A(register_addr[1]), .B(register_addr[0]), 
         .C(rw), .Z(n32017)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i260_2_lut_rep_400_3_lut.init = 16'hfefe;
    LUT4 n32472_bdd_2_lut (.A(n32472), .B(n1468[4]), .Z(n32473)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n32472_bdd_2_lut.init = 16'heeee;
    LUT4 n31984_bdd_4_lut_23773 (.A(n31984), .B(n32044), .C(n1468[0]), 
         .D(n1468[3]), .Z(n32472)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n31984_bdd_4_lut_23773.init = 16'hee0f;
    LUT4 i4532_2_lut_3_lut_4_lut_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(register_addr[2]), .D(n32032), .Z(n11158)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4532_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_43 (.A(databus[15]), .B(n5_adj_14), .C(n1468[13]), 
         .D(n29697), .Z(n27863)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_43.init = 16'hffec;
    LUT4 select_2107_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1468[4]), 
         .C(rx_data[7]), .D(n29971), .Z(n5_adj_14)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(register_addr[1]), .B(register_addr[0]), 
         .C(prev_select_adj_2), .D(rw), .Z(n4_adj_16)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23159_2_lut_rep_369_2_lut_3_lut_4_lut (.A(register_addr[1]), .B(register_addr[0]), 
         .C(register_addr[3]), .D(register_addr[2]), .Z(n31986)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23159_2_lut_rep_369_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i3566_2_lut_rep_440 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32057)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3566_2_lut_rep_440.init = 16'h8888;
    LUT4 mux_1537_i5_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[4]), 
         .D(n224[4]), .Z(n3899[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i14725_3_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(n9_adj_17), 
         .D(sendcount[2]), .Z(n19[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;
    defparam i14725_3_lut_4_lut.init = 16'h7f8f;
    LUT4 mux_1537_i16_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[15]), 
         .D(n224[15]), .Z(n3899[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 Select_4186_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[28] ), 
         .D(n33683), .Z(n3)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4186_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_44 (.A(databus[16]), .B(n5_adj_18), .C(n1468[13]), 
         .D(n29679), .Z(n27862)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_44.init = 16'hffec;
    LUT4 select_2107_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1468[4]), 
         .C(rx_data[0]), .D(n29984), .Z(n5_adj_18)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1537_i4_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[3]), 
         .D(n224[3]), .Z(n3899[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut (.A(n27768), .B(\control_reg[7] ), .C(n32088), .Z(n34)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut.init = 16'h0808;
    LUT4 i3569_2_lut_rep_442 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32059)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3569_2_lut_rep_442.init = 16'heeee;
    LUT4 i2_4_lut_adj_45 (.A(databus[17]), .B(n5_adj_19), .C(n1468[13]), 
         .D(n29698), .Z(n27852)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_45.init = 16'hffec;
    LUT4 select_2107_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1468[4]), 
         .C(rx_data[1]), .D(n29984), .Z(n5_adj_19)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_403_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n32020)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_403_3_lut.init = 16'h1e1e;
    LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.A(register_addr[0]), .B(n31933), 
         .C(n31991), .D(n29916), .Z(n13647)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_46.init = 16'hf4f0;
    LUT4 i2_4_lut_adj_47 (.A(databus[18]), .B(n5_adj_20), .C(n1468[13]), 
         .D(n29699), .Z(n27848)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_47.init = 16'hffec;
    LUT4 select_2107_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1468[4]), 
         .C(rx_data[2]), .D(n29984), .Z(n5_adj_20)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_48 (.A(databus[19]), .B(n5_adj_21), .C(n1468[13]), 
         .D(n29700), .Z(n27897)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_48.init = 16'hffec;
    LUT4 select_2107_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1468[4]), 
         .C(rx_data[3]), .D(n29984), .Z(n5_adj_21)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1537_i3_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[2]), 
         .D(n224[2]), .Z(n3899[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i3356_2_lut_rep_444 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32061)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i3356_2_lut_rep_444.init = 16'h9999;
    LUT4 i14793_3_lut_4_lut (.A(register_addr[0]), .B(n31933), .C(n32005), 
         .D(\register[2][3] ), .Z(n5980)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14793_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i2_4_lut_adj_49 (.A(databus[20]), .B(n5_adj_22), .C(n1468[13]), 
         .D(n29701), .Z(n27861)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_49.init = 16'hffec;
    LUT4 n12932_bdd_4_lut_23366_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n31115)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n12932_bdd_4_lut_23366_4_lut.init = 16'h6420;
    LUT4 select_2107_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1468[4]), 
         .C(rx_data[4]), .D(n29984), .Z(n5_adj_22)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_50 (.A(databus[21]), .B(n5_adj_23), .C(n1468[13]), 
         .D(n29702), .Z(n27847)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_50.init = 16'hffec;
    LUT4 i14726_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_adj_17), .Z(n19[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i14726_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 select_2107_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1468[4]), 
         .C(rx_data[5]), .D(n29984), .Z(n5_adj_23)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_51 (.A(databus[22]), .B(n5_adj_24), .C(n1468[13]), 
         .D(n29703), .Z(n27860)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_51.init = 16'hffec;
    LUT4 select_2107_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1468[4]), 
         .C(rx_data[6]), .D(n29984), .Z(n5_adj_24)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_52 (.A(databus[23]), .B(n5_adj_25), .C(n1468[13]), 
         .D(n29704), .Z(n27849)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_52.init = 16'hffec;
    LUT4 select_2107_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1468[4]), 
         .C(rx_data[7]), .D(n29984), .Z(n5_adj_25)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1537_i1_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[0]), 
         .D(n224[0]), .Z(n3899[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_53 (.A(databus[24]), .B(n5_adj_26), .C(n1468[13]), 
         .D(n29705), .Z(n27845)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_53.init = 16'hffec;
    LUT4 select_2107_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1468[4]), 
         .C(rx_data[0]), .D(n29983), .Z(n5_adj_26)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_54 (.A(databus[25]), .B(n5_adj_27), .C(n1468[13]), 
         .D(n29706), .Z(n27836)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_54.init = 16'hffec;
    LUT4 select_2107_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1468[4]), 
         .C(rx_data[1]), .D(n29983), .Z(n5_adj_27)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_55 (.A(databus[26]), .B(n5_adj_28), .C(n1468[13]), 
         .D(n29707), .Z(n27856)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_55.init = 16'hffec;
    LUT4 i1_2_lut_adj_56 (.A(n1468[16]), .B(n1468[19]), .Z(n2219)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_56.init = 16'heeee;
    LUT4 select_2107_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1468[4]), 
         .C(rx_data[2]), .D(n29983), .Z(n5_adj_28)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_57 (.A(databus[27]), .B(n5_adj_29), .C(n1468[13]), 
         .D(n29708), .Z(n27855)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_57.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_adj_58 (.A(rx_data[1]), .B(rx_data[4]), .C(rx_data[3]), 
         .Z(n13177)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_58.init = 16'h0808;
    LUT4 select_2107_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1468[4]), 
         .C(rx_data[3]), .D(n29983), .Z(n5_adj_29)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i2_3_lut_adj_59 (.A(n27787), .B(\control_reg[7]_adj_3 ), .C(n32088), 
         .Z(n32)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_59.init = 16'h0808;
    LUT4 i1_3_lut (.A(\select[4] ), .B(n33683), .C(prev_select_adj_4), 
         .Z(n29916)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut.init = 16'h0202;
    FD1P3IX send_491 (.D(n33682), .SP(n2219), .CD(n27886), .CK(debug_c_c), 
            .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 mux_1537_i10_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[9]), 
         .D(n224[9]), .Z(n3899[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_60 (.A(databus[28]), .B(n5_adj_32), .C(n1468[13]), 
         .D(n29709), .Z(n27822)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_60.init = 16'hffec;
    LUT4 select_2107_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1468[4]), 
         .C(rx_data[4]), .D(n29983), .Z(n5_adj_32)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_61 (.A(databus[29]), .B(n5_adj_33), .C(n1468[13]), 
         .D(n29682), .Z(n27824)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_61.init = 16'hffec;
    LUT4 n12932_bdd_2_lut_23376 (.A(sendcount[0]), .B(sendcount[3]), .Z(n31111)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n12932_bdd_2_lut_23376.init = 16'hbbbb;
    LUT4 select_2107_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1468[4]), 
         .C(rx_data[5]), .D(n29983), .Z(n5_adj_33)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut (.A(n1468[15]), .B(n7_adj_34), .C(n31118), .D(n30136), 
         .Z(n2738)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'h0020;
    LUT4 i14949_2_lut_rep_321_3_lut_4_lut (.A(register_addr[2]), .B(n32032), 
         .C(\select[4] ), .D(n13323), .Z(n31938)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14949_2_lut_rep_321_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_4189_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[27] ), 
         .D(n33683), .Z(n3_adj_5)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4189_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_62 (.A(register_addr[2]), .B(n32032), 
         .C(register_addr[1]), .D(n13323), .Z(n29798)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_62.init = 16'h0100;
    LUT4 mux_1537_i11_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[10]), 
         .D(n224[10]), .Z(n3899[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_320_3_lut_4_lut (.A(register_addr[2]), .B(n32032), 
         .C(register_addr[1]), .D(register_addr[5]), .Z(n31937)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_320_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_63 (.A(databus[30]), .B(n5_adj_36), .C(n1468[13]), 
         .D(n29680), .Z(n27842)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_63.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_64 (.A(register_addr[2]), .B(n32032), 
         .C(n32056), .D(n33680), .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_64.init = 16'hfffe;
    LUT4 select_2107_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1468[4]), 
         .C(rx_data[6]), .D(n29983), .Z(n5_adj_36)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_323_3_lut_4_lut (.A(register_addr[2]), .B(n32032), 
         .C(register_addr[1]), .D(n33680), .Z(n31940)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_323_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_316_3_lut_4_lut (.A(n32032), .B(n33680), .C(register_addr[1]), 
         .D(register_addr[2]), .Z(n31933)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_316_3_lut_4_lut.init = 16'h0010;
    LUT4 i23119_3_lut_4_lut (.A(n32032), .B(n33680), .C(register_addr[2]), 
         .D(n32056), .Z(n250_adj_6)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i23119_3_lut_4_lut.init = 16'h0111;
    LUT4 i1_3_lut_4_lut_rep_388 (.A(n32032), .B(n33680), .C(n32056), .D(register_addr[2]), 
         .Z(n32005)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_4_lut_rep_388.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_adj_65 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29984)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_65.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_66 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29983)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_66.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_461 (.A(\select[4] ), .B(register_addr[4]), .Z(n32078)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_461.init = 16'h8888;
    LUT4 i1_2_lut_rep_365_4_lut (.A(n167), .B(register_addr[3]), .C(n32034), 
         .D(n32090), .Z(n31982)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_365_4_lut.init = 16'h0002;
    LUT4 i2_3_lut_4_lut_adj_67 (.A(\select[4] ), .B(register_addr[4]), .C(n33683), 
         .D(prev_select_adj_2), .Z(n29904)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_67.init = 16'h0008;
    LUT4 i2_4_lut_adj_68 (.A(databus[31]), .B(n5_adj_38), .C(n1468[13]), 
         .D(n29710), .Z(n27838)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_68.init = 16'hffec;
    LUT4 select_2107_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1468[4]), 
         .C(rx_data[7]), .D(n29983), .Z(n5_adj_38)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n32046), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_adj_39)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_69 (.A(bufcount[0]), .B(n32046), .C(\buffer[0] [1]), 
         .D(rx_data[1]), .Z(n11_adj_40)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_69.init = 16'hf1e0;
    LUT4 i2_3_lut_4_lut_adj_70 (.A(register_addr[1]), .B(n31955), .C(n31972), 
         .D(n29904), .Z(n4071)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut_adj_70.init = 16'h0800;
    LUT4 i24_3_lut_4_lut_adj_71 (.A(bufcount[0]), .B(n32046), .C(\buffer[0] [2]), 
         .D(rx_data[2]), .Z(n11_adj_41)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_71.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_72 (.A(bufcount[0]), .B(n32046), .C(\buffer[0] [3]), 
         .D(rx_data[3]), .Z(n11_adj_42)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_72.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_73 (.A(bufcount[0]), .B(n32046), .C(rx_data[4]), 
         .D(\buffer[0] [4]), .Z(n11_adj_43)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_73.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_74 (.A(bufcount[0]), .B(n32046), .C(\buffer[0] [5]), 
         .D(rx_data[5]), .Z(n11_adj_44)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_74.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_75 (.A(bufcount[0]), .B(n32046), .C(rx_data[6]), 
         .D(\buffer[0] [6]), .Z(n11_adj_45)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_75.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_76 (.A(bufcount[0]), .B(n32046), .C(rx_data[7]), 
         .D(\buffer[0] [7]), .Z(n11_adj_46)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_76.init = 16'hfe10;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n32061), .B(n32020), .C(n4_adj_47), 
         .D(n32105), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n32061), .B(n32020), .C(n4_adj_48), 
         .D(n32108), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n32061), .B(n32020), .C(n4_adj_49), 
         .D(n32111), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n32061), .B(n32020), .C(n4_adj_50), 
         .D(n32117), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_1537_i12_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[11]), 
         .D(n224[11]), .Z(n3899[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i3312_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n31962), .C(n32018), 
         .D(bufcount[0]), .Z(n1864[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3312_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    LUT4 mux_1537_i13_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[12]), 
         .D(n224[12]), .Z(n3899[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_77 (.A(n1468[6]), .B(n1468[11]), .Z(n1921)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_77.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_78 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29972)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_78.init = 16'hfbfb;
    LUT4 i3_4_lut (.A(\buffer[0] [3]), .B(\buffer[0] [5]), .C(\buffer[0] [4]), 
         .D(\buffer[0] [6]), .Z(n12_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_79 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29971)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_79.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_80 (.A(n1468[3]), .B(n31984), .C(n1468[13]), 
         .Z(n14_c)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_80.init = 16'hf8f8;
    LUT4 i1_4_lut_adj_81 (.A(n1468[4]), .B(\buffer[0] [1]), .C(n11_adj_40), 
         .D(n14_c), .Z(n28826)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_81.init = 16'heca0;
    LUT4 i14734_2_lut_3_lut (.A(n1468[0]), .B(n1468[8]), .C(\select[2] ), 
         .Z(n16363)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14734_2_lut_3_lut.init = 16'h1010;
    LUT4 i14741_2_lut_3_lut (.A(n1468[0]), .B(n1468[8]), .C(\select[4] ), 
         .Z(n15376)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14741_2_lut_3_lut.init = 16'h1010;
    LUT4 i14745_2_lut_3_lut (.A(n1468[0]), .B(n1468[8]), .C(\select[3] ), 
         .Z(n15366)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14745_2_lut_3_lut.init = 16'h1010;
    LUT4 i14742_2_lut_3_lut (.A(n1468[0]), .B(n1468[8]), .C(\select[7] ), 
         .Z(n15372)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14742_2_lut_3_lut.init = 16'h1010;
    LUT4 i14738_2_lut_3_lut (.A(n1468[0]), .B(n1468[8]), .C(\select[1] ), 
         .Z(n16361)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14738_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_3_lut_4_lut_adj_82 (.A(n31983), .B(n29889), .C(prev_select_adj_4), 
         .D(n31991), .Z(n13708)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_82.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_adj_83 (.A(register_addr[5]), .B(n32003), .C(register_addr[1]), 
         .D(\select[4] ), .Z(n29883)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_83.init = 16'h2000;
    LUT4 i1_2_lut_4_lut_adj_84 (.A(register_addr[5]), .B(n32003), .C(register_addr[1]), 
         .D(register_addr[4]), .Z(n94)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_84.init = 16'h2000;
    LUT4 mux_1537_i17_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[16]), 
         .D(n224[16]), .Z(n3899[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_85 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [0]), 
         .Z(n29684)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_85.init = 16'h8080;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n32061), .B(n32020), .C(n4_adj_51), 
         .D(n32123), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n32061), .B(n32020), .C(n4_adj_52), 
         .D(n32120), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1468[4]), .B(n32045), .C(bufcount[0]), 
         .D(n31962), .Z(n27964)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hd222;
    LUT4 i1_4_lut_adj_86 (.A(n1468[4]), .B(\buffer[0] [2]), .C(n11_adj_41), 
         .D(n14_c), .Z(n28822)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_86.init = 16'heca0;
    LUT4 n31115_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n32059), .C(n32102), 
         .D(n31115), .Z(n31116)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n31115_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 mux_1537_i18_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[17]), 
         .D(n224[17]), .Z(n3899[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n32061), .B(n32020), .C(n4_adj_53), 
         .D(n32114), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_4_lut_adj_87 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][4] ), .Z(n29197)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_87.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_88 (.A(n32046), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n13275), .Z(n29673)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_88.init = 16'h0e00;
    LUT4 i23139_3_lut_4_lut (.A(n12_c), .B(\buffer[0] [2]), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n29981)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23139_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_4_lut_adj_89 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][5] ), .Z(n29211)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_89.init = 16'h0400;
    LUT4 i23153_3_lut_4_lut (.A(n12_c), .B(\buffer[0] [2]), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n29980)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23153_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_4_lut_adj_90 (.A(n1468[4]), .B(\buffer[0] [3]), .C(n11_adj_42), 
         .D(n14_c), .Z(n28836)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_90.init = 16'heca0;
    LUT4 i1_2_lut_4_lut_adj_91 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][6] ), .Z(n29213)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_91.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_92 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][7] ), .Z(n29207)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_92.init = 16'h0400;
    LUT4 i1_4_lut_adj_93 (.A(n1468[4]), .B(\buffer[0] [4]), .C(n11_adj_43), 
         .D(n14_c), .Z(n28858)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_93.init = 16'heca0;
    LUT4 i1_2_lut_4_lut_adj_94 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][8] ), .Z(n29199)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_94.init = 16'h0400;
    LUT4 i1_4_lut_adj_95 (.A(n1468[4]), .B(\buffer[0] [5]), .C(n11_adj_44), 
         .D(n14_c), .Z(n28814)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_95.init = 16'heca0;
    LUT4 i1_2_lut_4_lut_adj_96 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][9] ), .Z(n29215)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_96.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_97 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][10] ), .Z(n29189)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_97.init = 16'h0400;
    LUT4 i1_2_lut_rep_298_3_lut_4_lut (.A(register_addr[1]), .B(n31965), 
         .C(n29916), .D(register_addr[0]), .Z(n31915)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_298_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_4_lut_adj_98 (.A(n1468[4]), .B(\buffer[0] [6]), .C(n11_adj_45), 
         .D(n14_c), .Z(n28844)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_98.init = 16'heca0;
    LUT4 i1_4_lut_adj_99 (.A(n1468[4]), .B(\buffer[0] [7]), .C(n11_adj_46), 
         .D(n14_c), .Z(n28842)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_99.init = 16'heca0;
    LUT4 i1_4_lut_adj_100 (.A(n1468[4]), .B(\buffer[1] [0]), .C(n11_adj_54), 
         .D(n14_c), .Z(n28834)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_100.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_adj_101 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [1]), 
         .Z(n29686)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_101.init = 16'h8080;
    LUT4 i1_4_lut_adj_102 (.A(n32021), .B(debug_c_7), .C(n13275), .D(n8_adj_55), 
         .Z(n29014)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_102.init = 16'hdc50;
    LUT4 i1_4_lut_adj_103 (.A(n1468[4]), .B(\buffer[1] [1]), .C(n11_adj_56), 
         .D(n14_c), .Z(n28900)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_103.init = 16'heca0;
    LUT4 i14967_2_lut_rep_373_4_lut (.A(n32090), .B(register_addr[4]), .C(register_addr[5]), 
         .D(\select[3] ), .Z(n31990)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14967_2_lut_rep_373_4_lut.init = 16'h0400;
    LUT4 i1_3_lut_adj_104 (.A(n15_adj_57), .B(n1468[1]), .C(n1468[0]), 
         .Z(n8_adj_55)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut_adj_104.init = 16'hecec;
    LUT4 i1_2_lut_4_lut_adj_105 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][11] ), .Z(n29190)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_105.init = 16'h0400;
    LUT4 i15217_2_lut_rep_384_4_lut (.A(n32090), .B(register_addr[4]), .C(register_addr[5]), 
         .D(\select[3] ), .Z(n32001)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;
    defparam i15217_2_lut_rep_384_4_lut.init = 16'hfb00;
    LUT4 i3_4_lut_adj_106 (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), 
         .D(n29185), .Z(n15_adj_57)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i3_4_lut_adj_106.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_107 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [0]), 
         .Z(n29694)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_107.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_108 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][12] ), .Z(n29201)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_108.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_109 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][13] ), .Z(n29209)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_109.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_110 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][14] ), .Z(n29203)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_110.init = 16'h0400;
    LUT4 i3_4_lut_adj_111 (.A(n1468[3]), .B(n29663), .C(rx_data[2]), .D(n29835), 
         .Z(n13275)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_111.init = 16'h8000;
    LUT4 i2_4_lut_adj_112 (.A(escape), .B(n32042), .C(debug_c_7), .D(n13177), 
         .Z(n29663)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_4_lut_adj_112.init = 16'h1000;
    LUT4 i24_3_lut_4_lut_adj_113 (.A(bufcount[0]), .B(n32046), .C(\buffer[1] [0]), 
         .D(rx_data[0]), .Z(n11_adj_54)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_113.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_114 (.A(bufcount[0]), .B(n32046), .C(rx_data[1]), 
         .D(\buffer[1] [1]), .Z(n11_adj_56)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_114.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_adj_115 (.A(register_addr[1]), .B(n31965), 
         .C(n14372), .D(register_addr[0]), .Z(n9362)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_115.init = 16'h2000;
    LUT4 i1_4_lut_adj_116 (.A(n1468[4]), .B(\buffer[1] [2]), .C(n11_adj_58), 
         .D(n14_c), .Z(n28840)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_116.init = 16'heca0;
    LUT4 i1_4_lut_adj_117 (.A(sendcount[4]), .B(n1_c), .C(n6_adj_59), 
         .D(n12930), .Z(n9_adj_17)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_117.init = 16'hfeff;
    LUT4 i24_3_lut_4_lut_adj_118 (.A(bufcount[0]), .B(n32046), .C(\buffer[1] [2]), 
         .D(rx_data[2]), .Z(n11_adj_58)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_118.init = 16'hf2d0;
    LUT4 i1_2_lut_4_lut_adj_119 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][15] ), .Z(n29191)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_119.init = 16'h0400;
    LUT4 i24_3_lut_4_lut_adj_120 (.A(bufcount[0]), .B(n32046), .C(rx_data[3]), 
         .D(\buffer[1] [3]), .Z(n11_adj_60)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_120.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_121 (.A(bufcount[0]), .B(n32046), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_61)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_121.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_122 (.A(bufcount[0]), .B(n32046), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_62)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_122.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_123 (.A(bufcount[0]), .B(n32046), .C(rx_data[6]), 
         .D(\buffer[1] [6]), .Z(n11_adj_63)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_123.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_124 (.A(bufcount[0]), .B(n32046), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_64)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_124.init = 16'hf2d0;
    LUT4 i23113_3_lut_4_lut (.A(\buffer[0] [2]), .B(n12_c), .C(\buffer[0] [0]), 
         .D(\buffer[0] [1]), .Z(n28076)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23113_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_125 (.A(\buffer[0] [2]), .B(n12_c), .C(\buffer[0] [1]), 
         .Z(n29922)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i1_2_lut_3_lut_adj_125.init = 16'hefef;
    LUT4 i1_2_lut_4_lut_adj_126 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][16] ), .Z(n29193)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_126.init = 16'h0400;
    LUT4 i1_4_lut_adj_127 (.A(n1468[4]), .B(\buffer[1] [3]), .C(n11_adj_60), 
         .D(n14_c), .Z(n28884)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_127.init = 16'heca0;
    LUT4 i1_2_lut_rep_476 (.A(register_addr[4]), .B(register_addr[5]), .Z(n33680)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_476.init = 16'heeee;
    LUT4 i1_4_lut_adj_128 (.A(n1468[4]), .B(\buffer[1] [4]), .C(n11_adj_61), 
         .D(n14_c), .Z(n28850)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_128.init = 16'heca0;
    LUT4 equal_64_i1_4_lut (.A(sendcount[0]), .B(n22), .C(n12), .D(n8_adj_7), 
         .Z(n1_c)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_64_i1_4_lut.init = 16'h5556;
    LUT4 i1_2_lut_4_lut_adj_129 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][17] ), .Z(n29205)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_129.init = 16'h0400;
    LUT4 i1_2_lut_adj_130 (.A(rx_data[0]), .B(rx_data[5]), .Z(n29835)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_130.init = 16'h2222;
    LUT4 i2_4_lut_adj_131 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n32068), .Z(n6_adj_59)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_131.init = 16'he7de;
    LUT4 i1_4_lut_adj_132 (.A(n1468[4]), .B(\buffer[1] [5]), .C(n11_adj_62), 
         .D(n14_c), .Z(n28824)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_132.init = 16'heca0;
    LUT4 i1_4_lut_adj_133 (.A(n1468[4]), .B(debug_c_7), .C(n1468[2]), 
         .D(n29605), .Z(n28988)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_133.init = 16'heeea;
    LUT4 i1_4_lut_adj_134 (.A(n1468[4]), .B(\buffer[1] [6]), .C(n11_adj_63), 
         .D(n14_c), .Z(n28916)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_134.init = 16'heca0;
    LUT4 i1_4_lut_adj_135 (.A(n15_adj_57), .B(n1468[3]), .C(n1468[0]), 
         .D(n30106), .Z(n29605)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_135.init = 16'h50dc;
    LUT4 i22702_3_lut (.A(n13148), .B(escape), .C(n15_adj_57), .Z(n30106)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i22702_3_lut.init = 16'hecec;
    LUT4 reduce_or_463_i1_3_lut_4_lut (.A(n32021), .B(n13275), .C(\buffer[0] [7]), 
         .D(n1468[9]), .Z(n1573)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_463_i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_4_lut_adj_136 (.A(n1468[4]), .B(\buffer[1] [7]), .C(n11_adj_64), 
         .D(n14_c), .Z(n28818)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_136.init = 16'heca0;
    LUT4 i23171_3_lut (.A(debug_c_7), .B(n2), .C(n1468[3]), .Z(n29600)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i23171_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_387_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(register_addr[3]), .D(n32090), .Z(n32004)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_387_3_lut_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_137 (.A(escape), .B(n29835), .C(n31675), .D(n32042), 
         .Z(n2)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_137.init = 16'h0040;
    LUT4 mux_1537_i19_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[18]), 
         .D(n224[18]), .Z(n3899[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i14943_3_lut_4_lut (.A(n31971), .B(n1486), .C(n9_adj_17), .D(sendcount[0]), 
         .Z(n18[0])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i14943_3_lut_4_lut.init = 16'h0ddd;
    PFUMX i23358 (.BLUT(n31116), .ALUT(n31111), .C0(n5811), .Z(n31117));
    LUT4 i23212_2_lut_3_lut_4_lut (.A(register_addr[1]), .B(n31972), .C(register_addr[0]), 
         .D(register_addr[4]), .Z(n27946)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23212_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_rep_334_3_lut_4_lut (.A(register_addr[3]), .B(n32089), 
         .C(n29889), .D(n32090), .Z(n31951)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_334_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_1537_i14_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[13]), 
         .D(n224[13]), .Z(n3899[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX i8738 (.BLUT(n15368), .ALUT(n1864[1]), .C0(n1869), .Z(n15369));
    LUT4 i2_4_lut_adj_138 (.A(databus[0]), .B(n5_adj_67), .C(n1468[13]), 
         .D(n29684), .Z(n27934)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_138.init = 16'hffec;
    LUT4 select_2107_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1468[4]), 
         .C(rx_data[0]), .D(n29972), .Z(n5_adj_67)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 i3_4_lut_adj_139 (.A(n32003), .B(n167), .C(n33683), .D(register_addr[4]), 
         .Z(n52)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i3_4_lut_adj_139.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_adj_140 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][18] ), .Z(n29194)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_140.init = 16'h0400;
    PFUMX i8758 (.BLUT(n15388), .ALUT(n27964), .C0(n1869), .Z(n15389));
    LUT4 reduce_or_469_i1_3_lut (.A(busy), .B(n1468[13]), .C(n1480), .Z(n1579)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_469_i1_3_lut.init = 16'hdcdc;
    LUT4 i1_2_lut_rep_360_3_lut_4_lut (.A(register_addr[3]), .B(n32089), 
         .C(n32078), .D(n32090), .Z(n31977)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_360_3_lut_4_lut.init = 16'h0010;
    LUT4 i471_2_lut (.A(n5811), .B(n1486), .Z(n1580)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i471_2_lut.init = 16'h4444;
    LUT4 i2_4_lut_adj_141 (.A(databus[1]), .B(n5_adj_68), .C(n1468[13]), 
         .D(n29686), .Z(n27872)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_141.init = 16'hffec;
    LUT4 i248_2_lut_rep_417 (.A(register_addr[2]), .B(register_addr[4]), 
         .Z(n32034)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i248_2_lut_rep_417.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_142 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][19] ), .Z(n29196)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_142.init = 16'h0400;
    LUT4 select_2107_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1468[4]), 
         .C(rx_data[1]), .D(n29972), .Z(n5_adj_68)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_4_lut_adj_143 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][20] ), .Z(n29198)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_143.init = 16'h0400;
    LUT4 i2_4_lut_adj_144 (.A(databus[2]), .B(n5_adj_69), .C(n1468[13]), 
         .D(n29687), .Z(n27926)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_144.init = 16'hffec;
    LUT4 i1_2_lut_rep_472 (.A(register_addr[2]), .B(register_addr[5]), .Z(n32089)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_472.init = 16'heeee;
    LUT4 i1_2_lut_rep_416_3_lut (.A(register_addr[2]), .B(register_addr[5]), 
         .C(register_addr[3]), .Z(n32033)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_416_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_145 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][21] ), .Z(n29200)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_145.init = 16'h0400;
    LUT4 select_2107_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1468[4]), 
         .C(rx_data[2]), .D(n29972), .Z(n5_adj_69)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2107_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i2_3_lut_rep_391_4_lut (.A(register_addr[2]), .B(register_addr[4]), 
         .C(register_addr[3]), .D(n167), .Z(n32008)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_391_4_lut.init = 16'h0100;
    LUT4 i22700_2_lut_rep_366_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[5]), 
         .C(n32090), .D(register_addr[3]), .Z(n31983)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22700_2_lut_rep_366_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[5]), 
         .C(n29889), .D(register_addr[3]), .Z(n6_adj_70)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_473 (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .Z(n32090)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_473.init = 16'heeee;
    LUT4 i4400_3_lut (.A(n1468[16]), .B(n2738), .C(busy), .Z(n11026)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4400_3_lut.init = 16'hcece;
    LUT4 i5522_3_lut (.A(busy), .B(n1483), .C(n1468[16]), .Z(n12151)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5522_3_lut.init = 16'ha8a8;
    LUT4 i2_4_lut_adj_146 (.A(n38), .B(busy), .C(n31230), .D(n1483), 
         .Z(n28948)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_146.init = 16'hfbfa;
    LUT4 i1_4_lut_adj_147 (.A(n1468[15]), .B(n7_adj_34), .C(n31218), .D(n30136), 
         .Z(n38)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_147.init = 16'haaa8;
    LUT4 i1_2_lut_3_lut_adj_148 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [2]), 
         .Z(n29687)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_148.init = 16'h8080;
    LUT4 i2_3_lut_rep_395_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[5]), .D(register_addr[4]), .Z(n32012)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i2_3_lut_rep_395_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_4_lut_adj_149 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][22] ), .Z(n29202)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_149.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_150 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][23] ), .Z(n29204)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_150.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_adj_151 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [3]), 
         .Z(n29688)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_151.init = 16'h8080;
    LUT4 mux_1537_i20_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[19]), 
         .D(n224[19]), .Z(n3899[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1537_i21_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[20]), 
         .D(n224[20]), .Z(n3899[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1537_i22_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[21]), 
         .D(n224[21]), .Z(n3899[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 i4375_3_lut (.A(n1468[19]), .B(n1468[18]), .C(busy), .Z(n11000)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4375_3_lut.init = 16'hcece;
    LUT4 i5631_3_lut (.A(busy), .B(n1480), .C(n1468[19]), .Z(n12261)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5631_3_lut.init = 16'ha8a8;
    LUT4 i2_3_lut_rep_413_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[5]), .D(register_addr[4]), .Z(n32030)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_413_4_lut.init = 16'h0100;
    LUT4 i22636_2_lut_rep_415_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[3]), .Z(n32032)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22636_2_lut_rep_415_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_386_3_lut_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[2]), .D(register_addr[3]), .Z(n32003)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_386_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_152 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [4]), 
         .Z(n29691)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_152.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_153 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][24] ), .Z(n29206)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_153.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_adj_154 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [5]), 
         .Z(n29685)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_154.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_155 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][25] ), .Z(n29208)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_155.init = 16'h0400;
    LUT4 mux_1537_i23_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[22]), 
         .D(n224[22]), .Z(n3899[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_156 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][26] ), .Z(n29210)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_156.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_157 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][27] ), .Z(n29214)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_157.init = 16'h0400;
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_158 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [6]), 
         .Z(n29689)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_158.init = 16'h8080;
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2798), .CK(debug_c_c), 
            .Q(register_addr[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 mux_1537_i24_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[23]), 
         .D(n224[23]), .Z(n3899[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 i956_2_lut (.A(n1468[5]), .B(n31996), .Z(n2800)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i956_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_159 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4_adj_8)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_159.init = 16'h4444;
    LUT4 mux_1537_i25_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[24]), 
         .D(n224[24]), .Z(n3899[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_160 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][28] ), .Z(n29216)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_160.init = 16'h0400;
    LUT4 mux_1537_i26_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[25]), 
         .D(n224[25]), .Z(n3899[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_161 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][29] ), .Z(n29195)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_161.init = 16'h0400;
    LUT4 mux_1879_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n5811), 
         .Z(n5802[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1879_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_53)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 mux_1537_i27_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[26]), 
         .D(n224[26]), .Z(n3899[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_162 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][30] ), .Z(n29192)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_162.init = 16'h0400;
    LUT4 mux_1537_i28_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[27]), 
         .D(n224[27]), .Z(n3899[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1537_i29_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[28]), 
         .D(n224[28]), .Z(n3899[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_163 (.A(n32006), .B(register_addr[1]), .C(register_addr[0]), 
         .D(\register[2][31] ), .Z(n29212)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_163.init = 16'h0400;
    LUT4 i2_3_lut_rep_336 (.A(n29904), .B(register_addr[0]), .C(n31987), 
         .Z(n31953)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_3_lut_rep_336.init = 16'h2020;
    LUT4 mux_1537_i30_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[29]), 
         .D(n224[29]), .Z(n3899[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_164 (.A(n29904), .B(register_addr[0]), .C(n31987), 
         .D(n31991), .Z(n14094)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_164.init = 16'hff20;
    LUT4 mux_1537_i31_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[30]), 
         .D(n224[30]), .Z(n3899[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1537_i32_3_lut_4_lut (.A(n31928), .B(n31911), .C(databus[31]), 
         .D(n224[31]), .Z(n3899[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1537_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_293_3_lut_4_lut (.A(n31911), .B(n31970), .C(register_addr[1]), 
         .D(register_addr[0]), .Z(n31910)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_293_3_lut_4_lut.init = 16'h0080;
    LUT4 esc_data_2__bdd_4_lut (.A(esc_data[2]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[4]), .Z(n31118)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam esc_data_2__bdd_4_lut.init = 16'h4801;
    LUT4 i508_2_lut (.A(n1468[3]), .B(n1468[4]), .Z(n1869)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i508_2_lut.init = 16'heeee;
    FD1P3IX buffer_0___i2 (.D(n28826), .SP(n12818), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n28822), .SP(n12818), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n28836), .SP(n12818), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n28858), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n28814), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n28844), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n28842), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n28834), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n28900), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n28840), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n28884), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n28850), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n28824), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n28916), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n28818), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n27934), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n27872), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n27926), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n27931), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n27929), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i22 (.D(n27933), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    FD1P3IX buffer_0___i23 (.D(n27927), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n27937), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n27885), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n27928), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n27889), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n27930), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n27906), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n27851), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n27870), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n27863), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n27862), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n27852), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n27848), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n27897), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n27861), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n27847), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n27860), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n27849), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n27845), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n27836), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n27856), .SP(n14791), .CD(n31966), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n27855), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n27822), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n27824), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n27842), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n27838), .SP(n14791), .CD(n33689), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_165 (.A(n31911), .B(n31970), .C(register_addr[1]), 
         .D(register_addr[0]), .Z(n13710)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_165.init = 16'h0008;
    PFUMX i8742 (.BLUT(n15372), .ALUT(n29981), .C0(n1921), .Z(n15373));
    FD1S3IX state_FSM_i2 (.D(n29014), .CK(debug_c_c), .CD(n33689), .Q(n1468[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n28988), .CK(debug_c_c), .CD(n31966), .Q(n1468[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n12149), .CK(debug_c_c), .CD(n33689), .Q(n1468[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n29600), .CK(debug_c_c), .CD(n33689), .Q(n1468[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n29673), .CK(debug_c_c), .CD(n33689), .Q(n1468[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1468[5]), .CK(debug_c_c), .CD(n33689), .Q(n1468[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1468[6]), .CK(debug_c_c), .CD(n33689), .Q(n1468[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1468[7]), .CK(debug_c_c), .CD(n33689), .Q(n1468[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1468[8]), .CK(debug_c_c), .CD(n33689), 
            .Q(n1468[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1573), .CK(debug_c_c), .CD(n33689), .Q(n1468[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1468[10]), .CK(debug_c_c), .CD(n33689), 
            .Q(n1468[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1468[11]), .CK(debug_c_c), .CD(n33689), 
            .Q(n1468[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1468[12]), .CK(debug_c_c), .CD(n33689), 
            .Q(n1468[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1579), .CK(debug_c_c), .CD(n33689), .Q(n1486));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1580), .CK(debug_c_c), .CD(n33689), .Q(n1468[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n11026), .CK(debug_c_c), .CD(n33689), .Q(n1468[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n12151), .CK(debug_c_c), .CD(n33689), .Q(n1483));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n28948), .CK(debug_c_c), .CD(n33689), .Q(n1468[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n11000), .CK(debug_c_c), .CD(n33689), .Q(n1468[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i21 (.D(n12261), .CK(debug_c_c), .CD(n33689), .Q(n1480));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    LUT4 mux_1879_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n5811), 
         .Z(n5802[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1879_i3_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_52)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_adj_166 (.A(n1468[3]), .B(n31984), .C(\buffer[2] [7]), 
         .Z(n29681)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_166.init = 16'h8080;
    LUT4 i2_2_lut_adj_167 (.A(esc_data[7]), .B(esc_data[0]), .Z(n7_adj_34)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut_adj_167.init = 16'hbbbb;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_adj_51)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 mux_1879_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n5811), 
         .Z(n5802[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1879_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_168 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [1]), 
         .Z(n29690)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_168.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_169 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [2]), 
         .Z(n29693)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_169.init = 16'h8080;
    LUT4 i22732_2_lut (.A(esc_data[5]), .B(esc_data[6]), .Z(n30136)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22732_2_lut.init = 16'heeee;
    PFUMX i8746 (.BLUT(n15376), .ALUT(n29980), .C0(n1921), .Z(n15377));
    LUT4 mux_522_i4_3_lut (.A(n2738), .B(esc_data[3]), .C(n1468[18]), 
         .Z(n2210[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i4_3_lut.init = 16'hcaca;
    PFUMX i9731 (.BLUT(n16361), .ALUT(n28076), .C0(n1921), .Z(n16362));
    LUT4 Select_4192_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[26] ), 
         .D(n33683), .Z(n3_adj_9)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4192_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4195_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[25] ), 
         .D(n33683), .Z(n3_adj_10)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4195_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_522_i1_3_lut (.A(n2738), .B(esc_data[0]), .C(n1468[18]), 
         .Z(n2210[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i1_3_lut.init = 16'hcaca;
    LUT4 Select_4198_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[24] ), 
         .D(n33683), .Z(n3_adj_11)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4198_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_adj_170 (.A(register_addr[1]), .B(\steps_reg[5] ), .Z(n14)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_170.init = 16'h8888;
    LUT4 i1_2_lut_adj_171 (.A(register_addr[1]), .B(\steps_reg[6] ), .Z(n13)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_171.init = 16'h8888;
    LUT4 i1_2_lut_adj_172 (.A(register_addr[1]), .B(\steps_reg[3] ), .Z(n12_adj_12)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_172.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_173 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [3]), 
         .Z(n29692)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_173.init = 16'h8080;
    LUT4 Select_4201_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[23] ), 
         .D(rw), .Z(n3_adj_13)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4201_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i14618_2_lut (.A(sendcount[3]), .B(sendcount[0]), .Z(n9543[0])) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i14618_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_adj_174 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [4]), 
         .Z(n29695)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_174.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_175 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [5]), 
         .Z(n29696)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_175.init = 16'h8080;
    LUT4 Select_4204_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[22] ), 
         .D(rw), .Z(n3_adj_14)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4204_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_adj_176 (.A(register_addr[0]), .B(\control_reg[7]_adj_15 ), 
         .Z(n8494)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_176.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_177 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [6]), 
         .Z(n29683)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_177.init = 16'h8080;
    LUT4 Select_4207_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[21] ), 
         .D(rw), .Z(n3_adj_16)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4207_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_522_i2_3_lut (.A(n2738), .B(esc_data[1]), .C(n1468[18]), 
         .Z(n2210[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_178 (.A(n1468[3]), .B(n31984), .C(\buffer[3] [7]), 
         .Z(n29697)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_178.init = 16'h8080;
    LUT4 Select_4210_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[20] ), 
         .D(rw), .Z(n3_adj_17)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4210_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4213_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[19] ), 
         .D(rw), .Z(n3_adj_18)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4213_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4216_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[18] ), 
         .D(rw), .Z(n3_adj_19)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4216_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 \buffer_0[[0__bdd_4_lut_23661  (.A(\buffer[0] [0]), .B(n29922), 
         .C(n15366), .D(n1921), .Z(n31899)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam \buffer_0[[0__bdd_4_lut_23661 .init = 16'h22f0;
    LUT4 \buffer_0[[0__bdd_4_lut  (.A(\buffer[0] [0]), .B(n29922), .C(n16363), 
         .D(n1921), .Z(n31900)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam \buffer_0[[0__bdd_4_lut .init = 16'h11f0;
    LUT4 i1_2_lut_3_lut_adj_179 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [0]), 
         .Z(n29679)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_179.init = 16'h8080;
    LUT4 i3_4_lut_adj_180 (.A(n32017), .B(n6_adj_70), .C(prev_select_adj_4), 
         .D(n32090), .Z(n13642)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_4_lut_adj_180.init = 16'h0004;
    LUT4 i1_2_lut_adj_181 (.A(register_addr[0]), .B(\control_reg[7]_adj_20 ), 
         .Z(n8476)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_181.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_182 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [1]), 
         .Z(n29698)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_182.init = 16'h8080;
    LUT4 i14744_2_lut (.A(bufcount[1]), .B(n1468[0]), .Z(n15368)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14744_2_lut.init = 16'h2222;
    LUT4 Select_4219_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[17] ), 
         .D(rw), .Z(n3_adj_21)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4219_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i15703_3_lut_rep_343 (.A(n2738), .B(n31996), .C(n1468[18]), .Z(n31960)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15703_3_lut_rep_343.init = 16'hc8c8;
    LUT4 i23062_2_lut_3_lut (.A(n2738), .B(n31996), .C(n1468[18]), .Z(n16499)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i23062_2_lut_3_lut.init = 16'h0808;
    LUT4 Select_4222_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[16] ), 
         .D(rw), .Z(n3_adj_22)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4222_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4225_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[15] ), 
         .D(n33683), .Z(n3_adj_23)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4225_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4228_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[14] ), 
         .D(n33683), .Z(n3_adj_24)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4228_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_183 (.A(n32033), .B(n32078), .C(n32090), .D(n4_adj_16), 
         .Z(n13667)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_183.init = 16'h0004;
    LUT4 Select_4231_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[13] ), 
         .D(n33683), .Z(n3_adj_25)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4231_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_184 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [2]), 
         .Z(n29699)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_184.init = 16'h8080;
    LUT4 i2_4_lut_adj_185 (.A(n29883), .B(n31955), .C(n33683), .D(n4_adj_91), 
         .Z(n3984)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut_adj_185.init = 16'h0008;
    LUT4 i1_2_lut_adj_186 (.A(prev_select_adj_1), .B(register_addr[4]), 
         .Z(n4_adj_91)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_186.init = 16'heeee;
    LUT4 Select_4234_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[12] ), 
         .D(n33683), .Z(n3_adj_26)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4234_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_4_lut_adj_187 (.A(n5811), .B(n9543[0]), .C(n31996), .D(n1486), 
         .Z(n16497)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_187.init = 16'h8000;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n31960), .CD(n16499), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n31960), .CD(n16499), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n31960), .CD(n16499), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n31960), .CD(n16499), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n13608), .CD(n16497), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n13608), .CD(n16497), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n13608), .CD(n16497), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n13608), .CD(n16497), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=499, LSE_RLINE=509 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_50)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 Select_4237_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[11] ), 
         .D(n33683), .Z(n3_adj_27)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4237_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_49)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_188 (.A(n32008), .B(n32017), .C(prev_select_adj_1), 
         .D(n32090), .Z(n13693)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_188.init = 16'h0002;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_48)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_189 (.A(n29883), .B(rw), .C(n32052), .D(prev_select_adj_1), 
         .Z(n9139)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_4_lut_adj_189.init = 16'h0002;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_47)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_adj_190 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [3]), 
         .Z(n29700)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_190.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_191 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [4]), 
         .Z(n29701)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_191.init = 16'h8080;
    LUT4 i14740_2_lut (.A(bufcount[0]), .B(n1468[0]), .Z(n15388)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14740_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_adj_192 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [5]), 
         .Z(n29702)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_192.init = 16'h8080;
    LUT4 i1_2_lut_adj_193 (.A(register_addr[0]), .B(\control_reg[7] ), .Z(n1)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_193.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_194 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [6]), 
         .Z(n29703)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_194.init = 16'h8080;
    LUT4 i954_3_lut (.A(n1468[5]), .B(n31996), .C(n1468[10]), .Z(n2798)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i954_3_lut.init = 16'hc8c8;
    LUT4 i1_2_lut_3_lut_adj_195 (.A(n1468[3]), .B(n31984), .C(\buffer[4] [7]), 
         .Z(n29704)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_195.init = 16'h8080;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32095)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i2_3_lut_rep_325_4_lut (.A(register_addr[2]), .B(n32004), .C(rw), 
         .D(\select[4] ), .Z(n31942)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_rep_325_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_196 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [0]), 
         .Z(n29705)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_196.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_197 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [1]), 
         .Z(n29706)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_197.init = 16'h8080;
    LUT4 Select_4240_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[10] ), 
         .D(rw), .Z(n3_adj_28)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4240_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4243_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[9] ), 
         .D(n33683), .Z(n3_adj_29)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4243_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4246_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[8] ), 
         .D(n33683), .Z(n3_adj_30)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4246_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i5_3_lut (.A(n1468[9]), .B(n10), .C(n29997), .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_3_lut.init = 16'hfefe;
    LUT4 i4_4_lut (.A(n1468[15]), .B(n1483), .C(n1468[1]), .D(n32048), 
         .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_adj_198 (.A(n1468[19]), .B(n1468[3]), .C(n1468[11]), 
         .Z(n29997)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_adj_198.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_199 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [2]), 
         .Z(n29707)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_199.init = 16'h8080;
    LUT4 i1_4_lut_adj_200 (.A(n32047), .B(n1468[18]), .C(n8_adj_98), .D(n1468[6]), 
         .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_200.init = 16'hfffe;
    LUT4 i3_4_lut_adj_201 (.A(n1468[7]), .B(n1468[2]), .C(n29997), .D(n1468[10]), 
         .Z(n8_adj_98)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_201.init = 16'hfffe;
    LUT4 i2_3_lut_adj_202 (.A(n27766), .B(\control_reg[7]_adj_15 ), .C(n32088), 
         .Z(n32_adj_31)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_202.init = 16'h0808;
    LUT4 i4_4_lut_adj_203 (.A(n1468[4]), .B(n30007), .C(n1480), .D(n6), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_203.init = 16'hfffe;
    LUT4 i4_4_lut_adj_204 (.A(n1468[10]), .B(n8_adj_100), .C(n1468[13]), 
         .D(n30007), .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_204.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_205 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [3]), 
         .Z(n29708)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_205.init = 16'h8080;
    LUT4 i3_3_lut (.A(n1468[9]), .B(n1468[11]), .C(n1468[8]), .Z(n8_adj_100)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_3_lut.init = 16'hfefe;
    LUT4 i15701_3_lut_rep_354 (.A(n1468[13]), .B(n31996), .C(n1486), .Z(n31971)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15701_3_lut_rep_354.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_206 (.A(n1468[4]), .B(\buffer[0] [0]), .C(n11_adj_39), 
         .D(n14_c), .Z(n28838)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_206.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_adj_207 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [4]), 
         .Z(n29709)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_207.init = 16'h8080;
    LUT4 i23065_2_lut_rep_319_3_lut (.A(n1468[13]), .B(n31996), .C(n1486), 
         .Z(n31936)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i23065_2_lut_rep_319_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_adj_208 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [5]), 
         .Z(n29682)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_208.init = 16'h8080;
    LUT4 i1_3_lut_rep_304_4_lut (.A(register_addr[5]), .B(n32003), .C(n13700), 
         .D(register_addr[4]), .Z(n31921)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_rep_304_4_lut.init = 16'he0f0;
    LUT4 i23040_4_lut (.A(n7), .B(n30102), .C(n32044), .D(n1468[3]), 
         .Z(n12818)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i23040_4_lut.init = 16'h0544;
    LUT4 i22698_3_lut (.A(n1468[13]), .B(n1468[0]), .C(n1468[4]), .Z(n30102)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22698_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_209 (.A(register_addr[0]), .B(n31911), 
         .C(n31991), .D(register_addr[1]), .Z(n14661)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_209.init = 16'hf4f0;
    LUT4 i14724_4_lut (.A(sendcount[3]), .B(n9_adj_17), .C(sendcount[2]), 
         .D(n32057), .Z(n19[3])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(271[10:37])
    defparam i14724_4_lut.init = 16'h4888;
    LUT4 esc_data_1__bdd_4_lut (.A(esc_data[1]), .B(esc_data[3]), .C(esc_data[2]), 
         .D(esc_data[4]), .Z(n31218)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)))+!A (B+(C+(D)))) */ ;
    defparam esc_data_1__bdd_4_lut.init = 16'hd7fe;
    LUT4 i22778_4_lut (.A(rx_data[3]), .B(n32043), .C(rx_data[1]), .D(rx_data[4]), 
         .Z(n30186)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22778_4_lut.init = 16'hfffe;
    LUT4 i23132_2_lut_rep_305_3_lut_4_lut (.A(register_addr[5]), .B(n32003), 
         .C(register_addr[4]), .D(register_addr[1]), .Z(n31922)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i23132_2_lut_rep_305_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_adj_210 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [6]), 
         .Z(n29680)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_210.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_211 (.A(register_addr[5]), .B(n32003), 
         .C(register_addr[4]), .D(register_addr[1]), .Z(n96)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_211.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_212 (.A(n1468[3]), .B(n31984), .C(\buffer[5] [7]), 
         .Z(n29710)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_212.init = 16'h8080;
    LUT4 i15102_2_lut (.A(rx_data[2]), .B(rx_data[1]), .Z(n21696)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15102_2_lut.init = 16'heeee;
    PFUMX i23774 (.BLUT(n32474), .ALUT(n32473), .C0(bufcount[2]), .Z(n32475));
    LUT4 i1_4_lut_adj_213 (.A(n29715), .B(debug_c_7), .C(n1468[0]), .D(n1468[1]), 
         .Z(n13536)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_213.init = 16'hbbba;
    LUT4 n29714_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n31229)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n29714_bdd_4_lut.init = 16'h4001;
    LUT4 Select_4177_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[31] ), 
         .D(rw), .Z(n3_adj_32)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4177_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i3_4_lut_adj_214 (.A(sendcount[3]), .B(n32059), .C(sendcount[2]), 
         .D(n32041), .Z(n29715)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_214.init = 16'h0200;
    LUT4 Select_4183_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[29] ), 
         .D(rw), .Z(n3_adj_33)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4183_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_adj_215 (.A(register_addr[0]), .B(\control_reg[7]_adj_3 ), 
         .Z(n8485)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_215.init = 16'h4444;
    LUT4 i2_3_lut_4_lut_adj_216 (.A(n32078), .B(n31983), .C(prev_select_adj_2), 
         .D(n31991), .Z(n13700)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_216.init = 16'h0002;
    LUT4 Select_4180_i3_2_lut_3_lut_4_lut (.A(n32078), .B(n31983), .C(\read_value[30] ), 
         .D(rw), .Z(n3_adj_34)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4180_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n31986), .B(n32011), .C(n31990), .D(prev_select_adj_35), 
         .Z(n5)) /* synthesis lut_function=(!(A+!(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h5515;
    FD1P3AX rw_498_rep_477 (.D(n1468[10]), .SP(n2798), .CK(debug_c_c), 
            .Q(n33683));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_477.GSR = "ENABLED";
    PFUMX i23682 (.BLUT(n32121), .ALUT(n32122), .C0(sendcount[0]), .Z(n32123));
    PFUMX i23680 (.BLUT(n32118), .ALUT(n32119), .C0(sendcount[0]), .Z(n32120));
    PFUMX i23678 (.BLUT(n32115), .ALUT(n32116), .C0(sendcount[0]), .Z(n32117));
    PFUMX i23676 (.BLUT(n32112), .ALUT(n32113), .C0(sendcount[0]), .Z(n32114));
    PFUMX i23674 (.BLUT(n32109), .ALUT(n32110), .C0(sendcount[0]), .Z(n32111));
    PFUMX i23672 (.BLUT(n32106), .ALUT(n32107), .C0(sendcount[0]), .Z(n32108));
    PFUMX i23670 (.BLUT(n32103), .ALUT(n32104), .C0(sendcount[0]), .Z(n32105));
    LUT4 i23036_2_lut_2_lut (.A(n31996), .B(n12818), .Z(n14791)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i23036_2_lut_2_lut.init = 16'hdddd;
    PFUMX i23668 (.BLUT(n32100), .ALUT(n32101), .C0(sendcount[0]), .Z(n32102));
    PFUMX i23666 (.BLUT(n32097), .ALUT(n32098), .C0(n31962), .Z(n32099));
    PFUMX i23664 (.BLUT(n32094), .ALUT(n32095), .C0(sendcount[3]), .Z(n5811));
    LUT4 i2_3_lut_adj_217 (.A(n27769), .B(\control_reg[7]_adj_20 ), .C(n32088), 
         .Z(n32_adj_36)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_217.init = 16'h0808;
    \UARTTransmitter(baud_div=12)  uart_output (.n33689(n33689), .tx_data({tx_data}), 
            .n31996(n31996), .busy(busy), .\reset_count[14] (\reset_count[14] ), 
            .\reset_count[13] (\reset_count[13] ), .\reset_count[12] (\reset_count[12] ), 
            .n29900(n29900), .n31966(n31966), .send(send), .n10889(n10889), 
            .GND_net(GND_net), .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_c(debug_c_c), .n31996(n31996), 
            .rx_data({rx_data}), .n33689(n33689), .uart_rx_c(uart_rx_c), 
            .debug_c_7(debug_c_7), .n1497(n1468[3]), .n1498(n1468[2]), 
            .n12149(n12149), .n31966(n31966), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (n33689, tx_data, n31996, busy, 
            \reset_count[14] , \reset_count[13] , \reset_count[12] , n29900, 
            n31966, send, n10889, GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    output n33689;
    input [7:0]tx_data;
    output n31996;
    output busy;
    input \reset_count[14] ;
    input \reset_count[13] ;
    input \reset_count[12] ;
    input n29900;
    output n31966;
    input send;
    output n10889;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n31024;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9279, n17, n103, n2795, n31759, n31891, n31022, n31890, 
        n31514, n14695, n31023, n2, n30271, n7, n10, n29846, 
        n31958, n29847, n104, n30269, n30270, n29840, n4;
    
    FD1S3IX state__i0 (.D(n31024), .CK(bclk), .CD(n33689), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9279), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 i3_1_lut (.A(state[3]), .Z(n103)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i3_1_lut.init = 16'h5555;
    LUT4 n2794_bdd_4_lut (.A(n31996), .B(state[3]), .C(n2795), .D(state[2]), 
         .Z(n31759)) /* synthesis lut_function=(!((B (D)+!B !(C (D)))+!A)) */ ;
    defparam n2794_bdd_4_lut.init = 16'h2088;
    FD1P3IX busy_34 (.D(n103), .SP(n31891), .CD(n33689), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 i1_4_lut_rep_379 (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n29900), .Z(n31996)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i1_4_lut_rep_379.init = 16'heeea;
    LUT4 i15700_1_lut_rep_349_4_lut (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n29900), .Z(n31966)) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i15700_1_lut_rep_349_4_lut.init = 16'h1115;
    LUT4 state_1__bdd_2_lut (.A(state[0]), .B(state[3]), .Z(n31022)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 n31890_bdd_2_lut (.A(n31890), .B(state[2]), .Z(n31891)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n31890_bdd_2_lut.init = 16'h2222;
    LUT4 send_bdd_4_lut (.A(send), .B(state[3]), .C(state[1]), .D(state[0]), 
         .Z(n31514)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam send_bdd_4_lut.init = 16'h8001;
    LUT4 state_2__bdd_4_lut_23716 (.A(send), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n31890)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)))) */ ;
    defparam state_2__bdd_4_lut_23716.init = 16'hc002;
    LUT4 i23197_3_lut (.A(n31996), .B(n31514), .C(state[2]), .Z(n14695)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i23197_3_lut.init = 16'hf7f7;
    LUT4 state_1__bdd_4_lut_23457 (.A(state[1]), .B(state[0]), .C(send), 
         .D(state[3]), .Z(n31023)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;
    defparam state_1__bdd_4_lut_23457.init = 16'hb332;
    LUT4 i15700_1_lut_rep_483 (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n29900), .Z(n33689)) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i15700_1_lut_rep_483.init = 16'h1115;
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n30271), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15154_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15154_4_lut.init = 16'hfcee;
    FD1P3AX state__i3 (.D(n31759), .SP(n14695), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9279), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9279), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9279), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9279), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9279), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9279), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9279), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(n31996), .B(state[2]), .C(state[3]), .D(n2795), 
         .Z(n29846)) /* synthesis lut_function=(!((B (C+(D))+!B !(D))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2208;
    LUT4 i1_3_lut_rep_341 (.A(n31996), .B(state[2]), .C(state[3]), .Z(n31958)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut_rep_341.init = 16'h2a2a;
    LUT4 i1_3_lut (.A(state[1]), .B(n31958), .C(state[0]), .Z(n29847)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    FD1P3AX state__i2 (.D(n29846), .SP(n14695), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n29847), .SP(n14695), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 i22859_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n30269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22859_3_lut.init = 16'hcaca;
    LUT4 i22860_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n30270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22860_3_lut.init = 16'hcaca;
    PFUMX i22861 (.BLUT(n30269), .ALUT(n30270), .C0(state[1]), .Z(n30271));
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n33689), .CK(bclk), .Q(n10889)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    PFUMX i23313 (.BLUT(n31023), .ALUT(n31022), .C0(state[2]), .Z(n31024));
    LUT4 i951_2_lut (.A(state[0]), .B(state[1]), .Z(n2795)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i951_2_lut.init = 16'h8888;
    LUT4 i2_4_lut (.A(n29840), .B(state[2]), .C(n4), .D(n31996), .Z(n9279)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0200;
    LUT4 i1_2_lut (.A(send), .B(state[3]), .Z(n29840)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_adj_25 (.A(state[1]), .B(state[0]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_25.init = 16'heeee;
    \ClockDividerP(factor=12)  baud_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .bclk(bclk)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (GND_net, debug_c_c, bclk) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    output bclk;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    
    wire n27443, n8308, n27442;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27441, n27440, n27439, n27438, n27437, n27436, n27435, 
        n27434, n27433, n27432, n27431, n27430, n27429, n27428, 
        n30436, n49, n56, n50, n16539, n54, n46, n30204, n52, 
        n42, n48, n34, n27395;
    wire [31:0]n102;
    
    wire n27394, n27393, n27392, n27391, n27390, n27389, n27388, 
        n27387, n27386, n27385, n27384, n27383, n27382, n27381, 
        n27380;
    
    CCU2D sub_2056_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27443), .S0(n8308));
    defparam sub_2056_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2056_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2056_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2056_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27442), .COUT(n27443));
    defparam sub_2056_add_2_32.INIT0 = 16'h5555;
    defparam sub_2056_add_2_32.INIT1 = 16'h5555;
    defparam sub_2056_add_2_32.INJECT1_0 = "NO";
    defparam sub_2056_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27441), .COUT(n27442));
    defparam sub_2056_add_2_30.INIT0 = 16'h5555;
    defparam sub_2056_add_2_30.INIT1 = 16'h5555;
    defparam sub_2056_add_2_30.INJECT1_0 = "NO";
    defparam sub_2056_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27440), .COUT(n27441));
    defparam sub_2056_add_2_28.INIT0 = 16'h5555;
    defparam sub_2056_add_2_28.INIT1 = 16'h5555;
    defparam sub_2056_add_2_28.INJECT1_0 = "NO";
    defparam sub_2056_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27439), .COUT(n27440));
    defparam sub_2056_add_2_26.INIT0 = 16'h5555;
    defparam sub_2056_add_2_26.INIT1 = 16'h5555;
    defparam sub_2056_add_2_26.INJECT1_0 = "NO";
    defparam sub_2056_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27438), .COUT(n27439));
    defparam sub_2056_add_2_24.INIT0 = 16'h5555;
    defparam sub_2056_add_2_24.INIT1 = 16'h5555;
    defparam sub_2056_add_2_24.INJECT1_0 = "NO";
    defparam sub_2056_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27437), .COUT(n27438));
    defparam sub_2056_add_2_22.INIT0 = 16'h5555;
    defparam sub_2056_add_2_22.INIT1 = 16'h5555;
    defparam sub_2056_add_2_22.INJECT1_0 = "NO";
    defparam sub_2056_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27436), .COUT(n27437));
    defparam sub_2056_add_2_20.INIT0 = 16'h5555;
    defparam sub_2056_add_2_20.INIT1 = 16'h5555;
    defparam sub_2056_add_2_20.INJECT1_0 = "NO";
    defparam sub_2056_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27435), .COUT(n27436));
    defparam sub_2056_add_2_18.INIT0 = 16'h5555;
    defparam sub_2056_add_2_18.INIT1 = 16'h5555;
    defparam sub_2056_add_2_18.INJECT1_0 = "NO";
    defparam sub_2056_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27434), .COUT(n27435));
    defparam sub_2056_add_2_16.INIT0 = 16'h5555;
    defparam sub_2056_add_2_16.INIT1 = 16'h5555;
    defparam sub_2056_add_2_16.INJECT1_0 = "NO";
    defparam sub_2056_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27433), .COUT(n27434));
    defparam sub_2056_add_2_14.INIT0 = 16'h5555;
    defparam sub_2056_add_2_14.INIT1 = 16'h5555;
    defparam sub_2056_add_2_14.INJECT1_0 = "NO";
    defparam sub_2056_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27432), .COUT(n27433));
    defparam sub_2056_add_2_12.INIT0 = 16'h5555;
    defparam sub_2056_add_2_12.INIT1 = 16'h5555;
    defparam sub_2056_add_2_12.INJECT1_0 = "NO";
    defparam sub_2056_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27431), .COUT(n27432));
    defparam sub_2056_add_2_10.INIT0 = 16'h5555;
    defparam sub_2056_add_2_10.INIT1 = 16'h5555;
    defparam sub_2056_add_2_10.INJECT1_0 = "NO";
    defparam sub_2056_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27430), .COUT(n27431));
    defparam sub_2056_add_2_8.INIT0 = 16'h5555;
    defparam sub_2056_add_2_8.INIT1 = 16'h5555;
    defparam sub_2056_add_2_8.INJECT1_0 = "NO";
    defparam sub_2056_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27429), .COUT(n27430));
    defparam sub_2056_add_2_6.INIT0 = 16'h5555;
    defparam sub_2056_add_2_6.INIT1 = 16'h5555;
    defparam sub_2056_add_2_6.INJECT1_0 = "NO";
    defparam sub_2056_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27428), .COUT(n27429));
    defparam sub_2056_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2056_add_2_4.INIT1 = 16'h5555;
    defparam sub_2056_add_2_4.INJECT1_0 = "NO";
    defparam sub_2056_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2056_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27428));
    defparam sub_2056_add_2_2.INIT0 = 16'h0000;
    defparam sub_2056_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2056_add_2_2.INJECT1_0 = "NO";
    defparam sub_2056_add_2_2.INJECT1_1 = "NO";
    LUT4 i23126_4_lut (.A(n30436), .B(n49), .C(n56), .D(n50), .Z(n16539)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23126_4_lut.init = 16'h0002;
    LUT4 i23124_4_lut (.A(count[31]), .B(n54), .C(n46), .D(n30204), 
         .Z(n30436)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23124_4_lut.init = 16'h0100;
    LUT4 i19_4_lut (.A(count[24]), .B(count[27]), .C(count[4]), .D(count[30]), 
         .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(count[5]), .B(n52), .C(n42), .D(count[6]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i20_4_lut (.A(count[7]), .B(count[19]), .C(count[14]), .D(count[22]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(count[16]), .B(n48), .C(n34), .D(count[11]), 
         .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(count[28]), .B(count[2]), .C(count[18]), .D(count[8]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i22796_3_lut (.A(count[3]), .B(count[0]), .C(count[1]), .Z(n30204)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22796_3_lut.init = 16'h8080;
    LUT4 i18_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[21]), .B(count[25]), .Z(n34)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(count[15]), .B(count[29]), .C(count[23]), .D(count[13]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i12_2_lut (.A(count[10]), .B(count[20]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i12_2_lut.init = 16'heeee;
    CCU2D count_2641_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27395), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_33.INIT1 = 16'h0000;
    defparam count_2641_add_4_33.INJECT1_0 = "NO";
    defparam count_2641_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27394), .COUT(n27395), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_31.INJECT1_0 = "NO";
    defparam count_2641_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27393), .COUT(n27394), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_29.INJECT1_0 = "NO";
    defparam count_2641_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27392), .COUT(n27393), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_27.INJECT1_0 = "NO";
    defparam count_2641_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27391), .COUT(n27392), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_25.INJECT1_0 = "NO";
    defparam count_2641_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27390), .COUT(n27391), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_23.INJECT1_0 = "NO";
    defparam count_2641_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27389), .COUT(n27390), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_21.INJECT1_0 = "NO";
    defparam count_2641_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27388), .COUT(n27389), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_19.INJECT1_0 = "NO";
    defparam count_2641_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27387), .COUT(n27388), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_17.INJECT1_0 = "NO";
    defparam count_2641_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27386), .COUT(n27387), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_15.INJECT1_0 = "NO";
    defparam count_2641_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27385), .COUT(n27386), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_13.INJECT1_0 = "NO";
    defparam count_2641_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27384), .COUT(n27385), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_11.INJECT1_0 = "NO";
    defparam count_2641_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27383), .COUT(n27384), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_9.INJECT1_0 = "NO";
    defparam count_2641_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27382), .COUT(n27383), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_7.INJECT1_0 = "NO";
    defparam count_2641_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27381), .COUT(n27382), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_5.INJECT1_0 = "NO";
    defparam count_2641_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2641_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27380), .COUT(n27381), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2641_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2641_add_4_3.INJECT1_0 = "NO";
    defparam count_2641_add_4_3.INJECT1_1 = "NO";
    FD1S3IX count_2641__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i0.GSR = "ENABLED";
    CCU2D count_2641_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27380), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641_add_4_1.INIT0 = 16'hF000;
    defparam count_2641_add_4_1.INIT1 = 16'h0555;
    defparam count_2641_add_4_1.INJECT1_0 = "NO";
    defparam count_2641_add_4_1.INJECT1_1 = "NO";
    FD1S3AX clk_o_14 (.D(n8308), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2641__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i1.GSR = "ENABLED";
    FD1S3IX count_2641__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i2.GSR = "ENABLED";
    FD1S3IX count_2641__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i3.GSR = "ENABLED";
    FD1S3IX count_2641__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i4.GSR = "ENABLED";
    FD1S3IX count_2641__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i5.GSR = "ENABLED";
    FD1S3IX count_2641__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i6.GSR = "ENABLED";
    FD1S3IX count_2641__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i7.GSR = "ENABLED";
    FD1S3IX count_2641__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i8.GSR = "ENABLED";
    FD1S3IX count_2641__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i9.GSR = "ENABLED";
    FD1S3IX count_2641__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i10.GSR = "ENABLED";
    FD1S3IX count_2641__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i11.GSR = "ENABLED";
    FD1S3IX count_2641__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i12.GSR = "ENABLED";
    FD1S3IX count_2641__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i13.GSR = "ENABLED";
    FD1S3IX count_2641__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i14.GSR = "ENABLED";
    FD1S3IX count_2641__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i15.GSR = "ENABLED";
    FD1S3IX count_2641__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i16.GSR = "ENABLED";
    FD1S3IX count_2641__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i17.GSR = "ENABLED";
    FD1S3IX count_2641__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i18.GSR = "ENABLED";
    FD1S3IX count_2641__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i19.GSR = "ENABLED";
    FD1S3IX count_2641__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i20.GSR = "ENABLED";
    FD1S3IX count_2641__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i21.GSR = "ENABLED";
    FD1S3IX count_2641__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i22.GSR = "ENABLED";
    FD1S3IX count_2641__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i23.GSR = "ENABLED";
    FD1S3IX count_2641__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i24.GSR = "ENABLED";
    FD1S3IX count_2641__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i25.GSR = "ENABLED";
    FD1S3IX count_2641__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i26.GSR = "ENABLED";
    FD1S3IX count_2641__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i27.GSR = "ENABLED";
    FD1S3IX count_2641__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i28.GSR = "ENABLED";
    FD1S3IX count_2641__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i29.GSR = "ENABLED";
    FD1S3IX count_2641__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i30.GSR = "ENABLED";
    FD1S3IX count_2641__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16539), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2641__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_c, n31996, rx_data, n33689, 
            uart_rx_c, debug_c_7, n1497, n1498, n12149, n31966, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31996;
    output [7:0]rx_data;
    input n33689;
    input uart_rx_c;
    output debug_c_7;
    input n1497;
    input n1498;
    output n12149;
    input n31966;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n32035;
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n9227, n9229, n28912, baud_reset, n127, n32049, n32051, 
        n31985, bclk, n32050, n29988, n30118, n32, n31304, n31303, 
        n31317, n33631, n33632, n13334, n31318, n13, n9243, n10, 
        n28856, n29976;
    wire [7:0]n78;
    
    wire n9247, n32086, n9249, n130, n9251, n25408, n9253, n9255, 
        n13343, n19, n9257, n9259, n9261, n9263, n9265, n9267, 
        n9269, n24, n28, n31, n28372, n2, n10067;
    wire [5:0]n23;
    
    wire n16427, n29, n16428, n5, n21, n17, n28750, n31305, 
        n33633;
    
    LUT4 i3401_3_lut_rep_418 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n32035)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3401_3_lut_rep_418.init = 16'h8080;
    FD1P3AX rdata_i0_i0 (.D(n9227), .SP(n31996), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n9229), .SP(n31996), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n28912), .CK(debug_c_c), .CD(n33689), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n127), .CK(debug_c_c), .PD(n33689), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_432 (.A(state[1]), .B(state[4]), .Z(n32049)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_432.init = 16'heeee;
    LUT4 i1_2_lut_rep_368_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(uart_rx_c), 
         .D(n32051), .Z(n31985)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_368_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_433 (.A(state[1]), .B(bclk), .Z(n32050)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_rep_433.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut (.A(state[1]), .B(bclk), .C(state[3]), .Z(n29988)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i2_2_lut_rep_434 (.A(state[3]), .B(state[2]), .Z(n32051)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_rep_434.init = 16'heeee;
    LUT4 i22714_2_lut_3_lut (.A(state[3]), .B(state[2]), .C(uart_rx_c), 
         .Z(n30118)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22714_2_lut_3_lut.init = 16'hfefe;
    LUT4 n170_bdd_4_lut (.A(n31985), .B(state[1]), .C(n32), .D(state[5]), 
         .Z(n31304)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (D))) */ ;
    defparam n170_bdd_4_lut.init = 16'h00d5;
    LUT4 n170_bdd_2_lut (.A(state[1]), .B(bclk), .Z(n31303)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam n170_bdd_2_lut.init = 16'h9999;
    LUT4 n22036_bdd_4_lut (.A(uart_rx_c), .B(state[3]), .C(rdata[1]), 
         .D(state[2]), .Z(n31317)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)))) */ ;
    defparam n22036_bdd_4_lut.init = 16'hf0e2;
    LUT4 state_1__bdd_4_lut (.A(state[3]), .B(n32035), .C(state[4]), .D(bclk), 
         .Z(n33631)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;
    defparam state_1__bdd_4_lut.init = 16'hf078;
    LUT4 state_1__bdd_3_lut (.A(n32), .B(state[5]), .C(state[4]), .Z(n33632)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam state_1__bdd_3_lut.init = 16'h2020;
    LUT4 i1_4_lut (.A(n13334), .B(rdata[1]), .C(n31318), .D(n13), .Z(n9243)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_1 (.A(rdata[2]), .B(n13334), .C(n13), .D(n10), 
         .Z(n28856)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_1.init = 16'heca0;
    LUT4 i19_4_lut (.A(uart_rx_c), .B(rdata[2]), .C(n32050), .D(n29976), 
         .Z(n10)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i19_4_lut.init = 16'hccca;
    LUT4 i1_2_lut (.A(state[3]), .B(state[2]), .Z(n29976)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_2 (.A(n78[3]), .B(rdata[3]), .C(n13334), .D(n13), 
         .Z(n9247)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_2.init = 16'heca0;
    LUT4 i4366_4_lut (.A(uart_rx_c), .B(rdata[3]), .C(n32086), .D(n29976), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4366_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_3 (.A(n78[4]), .B(rdata[4]), .C(n13334), .D(n13), 
         .Z(n9249)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_3.init = 16'heca0;
    LUT4 i4364_4_lut (.A(uart_rx_c), .B(rdata[4]), .C(state[2]), .D(n29988), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4364_4_lut.init = 16'hccca;
    FD1S3IX drdy_51 (.D(n130), .CK(debug_c_c), .CD(n33689), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_4 (.A(n78[5]), .B(rdata[5]), .C(n13334), .D(n13), 
         .Z(n9251)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_4.init = 16'heca0;
    LUT4 i4362_4_lut (.A(uart_rx_c), .B(rdata[5]), .C(state[2]), .D(n25408), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4362_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_5 (.A(n78[6]), .B(rdata[6]), .C(n13334), .D(n13), 
         .Z(n9253)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_5.init = 16'heca0;
    LUT4 i4360_4_lut (.A(uart_rx_c), .B(rdata[6]), .C(state[2]), .D(n29988), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4360_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_6 (.A(n78[7]), .B(rdata[7]), .C(n13334), .D(n13), 
         .Z(n9255)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_6.init = 16'heca0;
    LUT4 i4358_4_lut (.A(rdata[7]), .B(uart_rx_c), .C(state[2]), .D(n25408), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4358_4_lut.init = 16'hcaaa;
    LUT4 i1_4_lut_adj_7 (.A(rdata[1]), .B(rx_data[1]), .C(n13343), .D(n19), 
         .Z(n9257)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_7.init = 16'heca0;
    LUT4 i1_4_lut_adj_8 (.A(rdata[2]), .B(rx_data[2]), .C(n13343), .D(n19), 
         .Z(n9259)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_8.init = 16'heca0;
    LUT4 i1_4_lut_adj_9 (.A(rdata[3]), .B(rx_data[3]), .C(n13343), .D(n19), 
         .Z(n9261)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_9.init = 16'heca0;
    LUT4 i1_4_lut_adj_10 (.A(rdata[4]), .B(rx_data[4]), .C(n13343), .D(n19), 
         .Z(n9263)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_10.init = 16'heca0;
    LUT4 i1_4_lut_adj_11 (.A(rdata[5]), .B(rx_data[5]), .C(n13343), .D(n19), 
         .Z(n9265)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_11.init = 16'heca0;
    LUT4 i1_4_lut_adj_12 (.A(rdata[6]), .B(rx_data[6]), .C(n13343), .D(n19), 
         .Z(n9267)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_12.init = 16'heca0;
    LUT4 i1_4_lut_adj_13 (.A(rdata[7]), .B(rx_data[7]), .C(n13343), .D(n19), 
         .Z(n9269)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_13.init = 16'heca0;
    LUT4 i45_4_lut (.A(n24), .B(n28), .C(state[5]), .D(n31), .Z(n28372)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i45_4_lut.init = 16'hfaca;
    LUT4 i3_3_lut_4_lut (.A(state[3]), .B(n32035), .C(bclk), .D(state[4]), 
         .Z(n2)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_4_lut_adj_14 (.A(state[4]), .B(state[0]), .C(state[1]), .D(n30118), 
         .Z(n28)) /* synthesis lut_function=(!(A+!(B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_14.init = 16'h4445;
    LUT4 i3415_2_lut_3_lut (.A(state[3]), .B(n32035), .C(state[4]), .Z(n10067)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3415_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_15 (.A(state[0]), .B(state[3]), .C(bclk), .D(n32035), 
         .Z(n31)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_15.init = 16'ha2aa;
    LUT4 mux_8_i4_3_lut_3_lut (.A(state[3]), .B(n32035), .C(bclk), .Z(n23[3])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam mux_8_i4_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i1_3_lut_4_lut (.A(state[0]), .B(n31985), .C(baud_reset), .D(n13343), 
         .Z(n127)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    defparam i1_3_lut_4_lut.init = 16'hffe0;
    LUT4 i9796_3_lut_3_lut (.A(state[3]), .B(n32035), .C(bclk), .Z(n16427)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i9796_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i1_3_lut_4_lut_adj_16 (.A(state[5]), .B(n32), .C(state[0]), .D(bclk), 
         .Z(n28912)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut_4_lut_adj_16.init = 16'hf400;
    LUT4 i2_3_lut_4_lut (.A(n32051), .B(n32049), .C(state[0]), .D(state[5]), 
         .Z(n13343)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i15436_2_lut_rep_469 (.A(bclk), .B(state[1]), .Z(n32086)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15436_2_lut_rep_469.init = 16'h8888;
    LUT4 rdata_1__bdd_3_lut_4_lut (.A(bclk), .B(state[1]), .C(n31317), 
         .D(rdata[1]), .Z(n31318)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam rdata_1__bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_17 (.A(bclk), .B(state[1]), .C(state[3]), 
         .Z(n25408)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_17.init = 16'h8080;
    LUT4 i1_3_lut (.A(debug_c_7), .B(n1497), .C(n1498), .Z(n12149)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut.init = 16'h5454;
    PFUMX i9797 (.BLUT(n29), .ALUT(n16427), .C0(state[0]), .Z(n16428));
    PFUMX i46 (.BLUT(n5), .ALUT(n2), .C0(state[0]), .Z(n24));
    PFUMX i32 (.BLUT(n21), .ALUT(n17), .C0(state[0]), .Z(n28750));
    FD1P3AX rdata_i0_i1 (.D(n9243), .SP(n31996), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n28856), .SP(n31996), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n9247), .SP(n31996), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n9249), .SP(n31996), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n9251), .SP(n31996), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n9253), .SP(n31996), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n9255), .SP(n31996), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n9257), .SP(n31996), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n9259), .SP(n31996), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n9261), .SP(n31996), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n9263), .SP(n31996), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n9265), .SP(n31996), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n9267), .SP(n31996), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n9269), .SP(n31996), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n31305), .CK(debug_c_c), .CD(n31966), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n28750), .CK(debug_c_c), .CD(n31966), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n16428), .CK(debug_c_c), .CD(n31966), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n33633), .CK(debug_c_c), .CD(n31966), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n28372), .CK(debug_c_c), .CD(n31966), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    PFUMX i24331 (.BLUT(n33632), .ALUT(n33631), .C0(state[0]), .Z(n33633));
    LUT4 i1_3_lut_4_lut_adj_18 (.A(state[0]), .B(n31985), .C(debug_c_7), 
         .D(n13343), .Z(n130)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    defparam i1_3_lut_4_lut_adj_18.init = 16'hffe0;
    LUT4 i20125_4_lut (.A(n23[3]), .B(state[5]), .C(n31985), .D(n32), 
         .Z(n29)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i20125_4_lut.init = 16'h2303;
    LUT4 i1_4_lut_adj_19 (.A(state[5]), .B(n32), .C(n10067), .D(bclk), 
         .Z(n5)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_19.init = 16'h4888;
    LUT4 i1_4_lut_adj_20 (.A(n78[0]), .B(rdata[0]), .C(n13334), .D(n13), 
         .Z(n9227)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_20.init = 16'heca0;
    LUT4 i4409_4_lut (.A(uart_rx_c), .B(rdata[0]), .C(n32051), .D(n32050), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4409_4_lut.init = 16'hccca;
    LUT4 i2_3_lut (.A(state[0]), .B(state[4]), .C(state[5]), .Z(n13334)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i2_3_lut_adj_21 (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_adj_21.init = 16'hefef;
    LUT4 i1_4_lut_adj_22 (.A(rdata[0]), .B(rx_data[0]), .C(n13343), .D(n19), 
         .Z(n9229)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_22.init = 16'heca0;
    LUT4 i4_4_lut (.A(n32051), .B(n32049), .C(state[5]), .D(state[0]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    LUT4 i1_4_lut_adj_23 (.A(state[4]), .B(state[2]), .C(state[3]), .D(state[1]), 
         .Z(n32)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_4_lut_adj_23.init = 16'heaaa;
    PFUMX i23421 (.BLUT(n31304), .ALUT(n31303), .C0(state[0]), .Z(n31305));
    LUT4 i1_4_lut_adj_24 (.A(state[5]), .B(state[2]), .C(n31985), .D(n32), 
         .Z(n21)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_24.init = 16'h4505;
    LUT4 i33_3_lut (.A(state[1]), .B(state[2]), .C(bclk), .Z(n17)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i33_3_lut.init = 16'hc6c6;
    \ClockDividerP(factor=12)_U0  baud_gen (.GND_net(GND_net), .bclk(bclk), 
            .debug_c_c(debug_c_c), .baud_reset(baud_reset)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (GND_net, bclk, debug_c_c, baud_reset) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output bclk;
    input debug_c_c;
    input baud_reset;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27459, n8273, n27458;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27457, n27456, n27455, n27454, n27453, n27452, n27451, 
        n27450, n27449, n27448, n27447, n27446, n27445, n27444, 
        n2950;
    wire [31:0]n134;
    
    wire n55, n27603, n56, n52, n44, n35, n54, n48, n36, n46, 
        n32, n50, n40, n27379, n27378, n27377, n27376, n27375, 
        n27374, n27373, n27372, n27371, n27370, n27369, n27368, 
        n27367, n27366, n27365, n27364;
    
    CCU2D sub_2054_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27459), .S0(n8273));
    defparam sub_2054_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2054_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2054_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2054_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27458), .COUT(n27459));
    defparam sub_2054_add_2_32.INIT0 = 16'h5555;
    defparam sub_2054_add_2_32.INIT1 = 16'h5555;
    defparam sub_2054_add_2_32.INJECT1_0 = "NO";
    defparam sub_2054_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27457), .COUT(n27458));
    defparam sub_2054_add_2_30.INIT0 = 16'h5555;
    defparam sub_2054_add_2_30.INIT1 = 16'h5555;
    defparam sub_2054_add_2_30.INJECT1_0 = "NO";
    defparam sub_2054_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27456), .COUT(n27457));
    defparam sub_2054_add_2_28.INIT0 = 16'h5555;
    defparam sub_2054_add_2_28.INIT1 = 16'h5555;
    defparam sub_2054_add_2_28.INJECT1_0 = "NO";
    defparam sub_2054_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27455), .COUT(n27456));
    defparam sub_2054_add_2_26.INIT0 = 16'h5555;
    defparam sub_2054_add_2_26.INIT1 = 16'h5555;
    defparam sub_2054_add_2_26.INJECT1_0 = "NO";
    defparam sub_2054_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27454), .COUT(n27455));
    defparam sub_2054_add_2_24.INIT0 = 16'h5555;
    defparam sub_2054_add_2_24.INIT1 = 16'h5555;
    defparam sub_2054_add_2_24.INJECT1_0 = "NO";
    defparam sub_2054_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27453), .COUT(n27454));
    defparam sub_2054_add_2_22.INIT0 = 16'h5555;
    defparam sub_2054_add_2_22.INIT1 = 16'h5555;
    defparam sub_2054_add_2_22.INJECT1_0 = "NO";
    defparam sub_2054_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27452), .COUT(n27453));
    defparam sub_2054_add_2_20.INIT0 = 16'h5555;
    defparam sub_2054_add_2_20.INIT1 = 16'h5555;
    defparam sub_2054_add_2_20.INJECT1_0 = "NO";
    defparam sub_2054_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27451), .COUT(n27452));
    defparam sub_2054_add_2_18.INIT0 = 16'h5555;
    defparam sub_2054_add_2_18.INIT1 = 16'h5555;
    defparam sub_2054_add_2_18.INJECT1_0 = "NO";
    defparam sub_2054_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27450), .COUT(n27451));
    defparam sub_2054_add_2_16.INIT0 = 16'h5555;
    defparam sub_2054_add_2_16.INIT1 = 16'h5555;
    defparam sub_2054_add_2_16.INJECT1_0 = "NO";
    defparam sub_2054_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27449), .COUT(n27450));
    defparam sub_2054_add_2_14.INIT0 = 16'h5555;
    defparam sub_2054_add_2_14.INIT1 = 16'h5555;
    defparam sub_2054_add_2_14.INJECT1_0 = "NO";
    defparam sub_2054_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27448), .COUT(n27449));
    defparam sub_2054_add_2_12.INIT0 = 16'h5555;
    defparam sub_2054_add_2_12.INIT1 = 16'h5555;
    defparam sub_2054_add_2_12.INJECT1_0 = "NO";
    defparam sub_2054_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27447), .COUT(n27448));
    defparam sub_2054_add_2_10.INIT0 = 16'h5555;
    defparam sub_2054_add_2_10.INIT1 = 16'h5555;
    defparam sub_2054_add_2_10.INJECT1_0 = "NO";
    defparam sub_2054_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27446), .COUT(n27447));
    defparam sub_2054_add_2_8.INIT0 = 16'h5555;
    defparam sub_2054_add_2_8.INIT1 = 16'h5555;
    defparam sub_2054_add_2_8.INJECT1_0 = "NO";
    defparam sub_2054_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27445), .COUT(n27446));
    defparam sub_2054_add_2_6.INIT0 = 16'h5555;
    defparam sub_2054_add_2_6.INIT1 = 16'h5555;
    defparam sub_2054_add_2_6.INJECT1_0 = "NO";
    defparam sub_2054_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27444), .COUT(n27445));
    defparam sub_2054_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2054_add_2_4.INIT1 = 16'h5555;
    defparam sub_2054_add_2_4.INJECT1_0 = "NO";
    defparam sub_2054_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27444));
    defparam sub_2054_add_2_2.INIT0 = 16'h0000;
    defparam sub_2054_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2054_add_2_2.INJECT1_0 = "NO";
    defparam sub_2054_add_2_2.INJECT1_1 = "NO";
    FD1S3IX clk_o_14 (.D(n8273), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2640__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2950), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i0.GSR = "ENABLED";
    LUT4 i1106_4_lut (.A(n55), .B(baud_reset), .C(n27603), .D(n56), 
         .Z(n2950)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i1106_4_lut.init = 16'hccdc;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(count[1]), .B(count[3]), .C(count[0]), .Z(n27603)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_2_lut.init = 16'heeee;
    CCU2D count_2640_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27379), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_33.INIT1 = 16'h0000;
    defparam count_2640_add_4_33.INJECT1_0 = "NO";
    defparam count_2640_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27378), .COUT(n27379), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_31.INJECT1_0 = "NO";
    defparam count_2640_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27377), .COUT(n27378), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_29.INJECT1_0 = "NO";
    defparam count_2640_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27376), .COUT(n27377), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_27.INJECT1_0 = "NO";
    defparam count_2640_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27375), .COUT(n27376), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_25.INJECT1_0 = "NO";
    defparam count_2640_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27374), .COUT(n27375), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_23.INJECT1_0 = "NO";
    defparam count_2640_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27373), .COUT(n27374), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_21.INJECT1_0 = "NO";
    defparam count_2640_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27372), .COUT(n27373), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_19.INJECT1_0 = "NO";
    defparam count_2640_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27371), .COUT(n27372), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_17.INJECT1_0 = "NO";
    defparam count_2640_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27370), .COUT(n27371), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_15.INJECT1_0 = "NO";
    defparam count_2640_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27369), .COUT(n27370), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_13.INJECT1_0 = "NO";
    defparam count_2640_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27368), .COUT(n27369), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_11.INJECT1_0 = "NO";
    defparam count_2640_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27367), .COUT(n27368), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_9.INJECT1_0 = "NO";
    defparam count_2640_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27366), .COUT(n27367), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_7.INJECT1_0 = "NO";
    defparam count_2640_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27365), .COUT(n27366), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_5.INJECT1_0 = "NO";
    defparam count_2640_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27364), .COUT(n27365), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2640_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2640_add_4_3.INJECT1_0 = "NO";
    defparam count_2640_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2640_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27364), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640_add_4_1.INIT0 = 16'hF000;
    defparam count_2640_add_4_1.INIT1 = 16'h0555;
    defparam count_2640_add_4_1.INJECT1_0 = "NO";
    defparam count_2640_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2640__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2950), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i1.GSR = "ENABLED";
    FD1S3IX count_2640__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2950), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i2.GSR = "ENABLED";
    FD1S3IX count_2640__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2950), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i3.GSR = "ENABLED";
    FD1S3IX count_2640__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2950), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i4.GSR = "ENABLED";
    FD1S3IX count_2640__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2950), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i5.GSR = "ENABLED";
    FD1S3IX count_2640__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2950), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i6.GSR = "ENABLED";
    FD1S3IX count_2640__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2950), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i7.GSR = "ENABLED";
    FD1S3IX count_2640__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2950), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i8.GSR = "ENABLED";
    FD1S3IX count_2640__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2950), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i9.GSR = "ENABLED";
    FD1S3IX count_2640__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i10.GSR = "ENABLED";
    FD1S3IX count_2640__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i11.GSR = "ENABLED";
    FD1S3IX count_2640__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i12.GSR = "ENABLED";
    FD1S3IX count_2640__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i13.GSR = "ENABLED";
    FD1S3IX count_2640__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i14.GSR = "ENABLED";
    FD1S3IX count_2640__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i15.GSR = "ENABLED";
    FD1S3IX count_2640__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i16.GSR = "ENABLED";
    FD1S3IX count_2640__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i17.GSR = "ENABLED";
    FD1S3IX count_2640__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i18.GSR = "ENABLED";
    FD1S3IX count_2640__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i19.GSR = "ENABLED";
    FD1S3IX count_2640__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i20.GSR = "ENABLED";
    FD1S3IX count_2640__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i21.GSR = "ENABLED";
    FD1S3IX count_2640__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i22.GSR = "ENABLED";
    FD1S3IX count_2640__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i23.GSR = "ENABLED";
    FD1S3IX count_2640__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i24.GSR = "ENABLED";
    FD1S3IX count_2640__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i25.GSR = "ENABLED";
    FD1S3IX count_2640__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i26.GSR = "ENABLED";
    FD1S3IX count_2640__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i27.GSR = "ENABLED";
    FD1S3IX count_2640__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i28.GSR = "ENABLED";
    FD1S3IX count_2640__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i29.GSR = "ENABLED";
    FD1S3IX count_2640__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i30.GSR = "ENABLED";
    FD1S3IX count_2640__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2950), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2640__i31.GSR = "ENABLED";
    
endmodule
