// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Thu Apr  7 01:28:40 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    output expansion4 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire n31780 /* synthesis SET_AS_NETWORK=n31780 */ ;
    wire n33445 /* synthesis nomerge= */ ;
    wire n31762 /* synthesis SET_AS_NETWORK=n31762 */ ;
    
    wire GND_net, VCC_net, n10608_c, n10607, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, signal_light_c, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
        encoder_la_c, encoder_lb_c, encoder_li_c, rc_ch1_c, rc_ch2_c, 
        rc_ch3_c, rc_ch4_c, rc_ch7_c, rc_ch8_c, motor_pwm_l_c, xbee_pause_c, 
        debug_c_7, debug_c_5, debug_c_4, debug_c_3, debug_c_2;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire rw, n14124, n27915, n24;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    wire [4:0]arm_select;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(523[12:22])
    
    wire clk_10Hz, n1, n34, n22093, n21, n30191, n14084, n31724, 
        n14194, n31722, n5, n22, n2, n5_adj_570, n20991, n20993, 
        n31695, n31694;
    wire [7:0]n8242;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n27902, n27385, n27384, n27383, n27382, n14022, n27381, 
        n22_adj_571, n27380, n32, n27379, n4, n6;
    wire [31:0]n1294;
    
    wire n27918, n14187, n14186, n14183, n14182, n5613, n8110, 
        n24311, n14176, n29, n30218, n14172, n32_adj_572, n30195, 
        n2669, n32_adj_573, n31720, n3, n3786;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[12:21])
    
    wire prev_select, n46, n31719, n24417;
    wire [7:0]\register[1]_adj_855 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]\register[0]_adj_856 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [2:0]read_size_adj_858;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(93[12:21])
    
    wire n30186, n30216, n29452, n29823, n27924, n27884, n2658, 
        n29694, n30197, n33448, n241, n8885;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched, prev_limit_latched, step_clk, prev_step_clk;
    wire [31:0]read_value_adj_864;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_865;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_609, n29853, n29850, n106, n185, n191;
    wire [31:0]n580;
    
    wire n3970;
    wire [7:0]control_reg_adj_873;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_874;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_875;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire int_step, step_clk_adj_611, prev_step_clk_adj_612;
    wire [31:0]read_value_adj_876;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_877;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_647, n3_adj_648, n27910, n30205, n5_adj_649, 
        n27905, n31718, n13779;
    wire [7:0]control_reg_adj_913;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire step_clk_adj_651, prev_step_clk_adj_652;
    wire [31:0]read_value_adj_916;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_917;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_687, n8940, n27893, n13757, n31717, n30184, 
        n8;
    wire [7:0]control_reg_adj_953;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]read_value_adj_956;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_957;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_723, n28025;
    wire [31:0]n99_adj_1259;
    wire [7:0]n571_adj_974;
    
    wire n6_adj_724, n31716, n21959;
    wire [31:0]read_value_adj_996;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[13:23])
    wire [2:0]read_size_adj_997;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(67[12:21])
    
    wire n47_adj_759;
    wire [2:0]n249;
    wire [31:0]read_value_adj_1005;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[13:23])
    wire [2:0]read_size_adj_1006;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(67[12:21])
    
    wire n28845, n2_adj_763, n31715, n1_adj_764, n3700, n30182, 
        n13719, n4_adj_765, n14252, n27707, n13671, n13606, n13568, 
        n30152, n28937, n29930, n9, n14, n10, n9_adj_766, n31713, 
        n6_adj_767, n3_adj_768, n2_adj_769, n5_adj_770, n8_adj_771;
    wire [14:0]n66_adj_1391;
    
    wire n8_adj_772, n2_adj_773, n5_adj_774, n6_adj_775, n2_adj_776, 
        n8_adj_777, n3_adj_778, n2_adj_779, n5_adj_780, n8_adj_781, 
        n2_adj_782, n5_adj_783, n8_adj_784, n3_adj_785, n3_adj_786, 
        n6_adj_787, n6_adj_788, n3_adj_789, n3_adj_790, n6_adj_791, 
        n6_adj_792, n6_adj_793, n3_adj_794, n6_adj_795, n3_adj_796, 
        n6_adj_797, n3_adj_798, n3_adj_799, n3_adj_800, n6_adj_801, 
        n6_adj_802, n3_adj_803, n6_adj_804, n3_adj_805, n6_adj_806, 
        n3_adj_807, n6_adj_808, n3_adj_809, n6_adj_810, n3_adj_811, 
        n6_adj_812, n3_adj_813, n6_adj_814, n3_adj_815, n33447, n31712, 
        n6_adj_816, n31711, n3_adj_817, n31708, n6_adj_818, n31707, 
        n31705, n31703, n31702, n6_adj_819, n3_adj_820, n6_adj_821, 
        n3_adj_822, n8_adj_823, n31701;
    wire [3:0]n7447;
    
    wire n31700, n12, n6_adj_824;
    wire [7:0]n8260;
    
    wire n30160;
    wire [7:0]n8251;
    
    wire n9_adj_825, n21892, n27937;
    wire [31:0]n6558;
    
    wire n30, n31867, n5_adj_826, n2_adj_827, n31699;
    wire [3:0]state_adj_1040;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    
    wire select_clk;
    wire [31:0]n15;
    wire [31:0]n59;
    
    wire n31841;
    wire [31:0]n99_adj_1262;
    
    wire n31832, n33457, n31237, n31827, n29738, n31818, n13476, 
        n21729, n33455, n31798, n9093, n31, n19, n31797, n31796, 
        n3883, n6_adj_829, n20980, n13, n33453, n24690, n20982, 
        n33452, n20983, n14_adj_830, n9089, n31785;
    wire [31:0]n4137;
    
    wire n31784, n31783, n24720, n24729, n33451, n31779, n24748, 
        n31698, n27912, n33450, n29552, n31774, n29370, n3_adj_831, 
        n33449, n78_adj_832, n89_adj_833, n27933, n17753, n17748, 
        n17745, n17735, n7485, n29966, n14424, n31763, n29590, 
        n9848, n31759, n16046, n16045, n33446, n31751;
    wire [3:0]state_adj_1182;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n31746, n30189, n31741, n31739, n12795, n31733, n31732, 
        n31727, n10675, n55;
    
    VHI i2 (.Z(VCC_net));
    GlobalControlPeripheral global_control (.\register[2] ({Open_0, Open_1, 
            Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, 
            Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
            Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, 
            Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, 
            Open_27, Open_28, Open_29, Open_30, \register[2] [0]}), 
            .debug_c_c(debug_c_c), .n33450(n33450), .read_size({read_size}), 
            .n14022(n14022), .n24748(n24748), .prev_select(prev_select), 
            .\select[1] (select[1]), .n33449(n33449), .n33446(n33446), 
            .n46(n46), .read_value({read_value}), .n28937(n28937), .GND_net(GND_net), 
            .n33448(n33448), .\databus[1] (databus[1]), .\register_addr[1] (register_addr[1]), 
            .n31739(n31739), .\register_addr[0] (register_addr[0]), .n27707(n27707), 
            .n31827(n31827), .n31702(n31702), .rw(rw), .n33447(n33447), 
            .n29823(n29823), .n24729(n24729), .n31720(n31720), .n31832(n31832), 
            .\control_reg[7] (control_reg_adj_873[7]), .n27893(n27893), 
            .n32(n32_adj_573), .\control_reg[7]_adj_301 (control_reg_adj_953[7]), 
            .n27905(n27905), .n32_adj_302(n32_adj_572), .n21959(n21959), 
            .\register[1][1] (\register[1]_adj_855 [1]), .n31796(n31796), 
            .signal_light_c(signal_light_c), .\control_reg[7]_adj_303 (control_reg_adj_913[7]), 
            .n27902(n27902), .n32_adj_304(n32), .\control_reg[7]_adj_305 (control_reg[7]), 
            .n27910(n27910), .n34(n34), .n21892(n21892), .\register[0][1] (\register[0]_adj_856 [1]), 
            .n31797(n31797), .\register[0][7] (\register[0]_adj_856 [7]), 
            .n31798(n31798), .n21729(n21729), .n31(n31), .\state[0] (state_adj_1040[0]), 
            .n19(n19), .\register_addr[2] (register_addr[2]), .n29738(n29738), 
            .n21(n21), .n31779(n31779), .\register_addr[5] (register_addr[5]), 
            .\register_addr[4] (register_addr[4]), .xbee_pause_c(xbee_pause_c), 
            .n16046(n16046), .n16045(n16045), .n31718(n31718), .n29452(n29452)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(495[45] 505[74])
    LUT4 i14620_3_lut (.A(Stepper_Y_Dir_c), .B(div_factor_reg_adj_874[5]), 
         .C(register_addr[1]), .Z(n20991)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i14620_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(state_adj_1182[2]), .B(n31237), .C(n33447), .Z(n14424)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    PFUMX i14622 (.BLUT(n20991), .ALUT(n14_adj_830), .C0(register_addr[0]), 
          .Z(n20993));
    LUT4 i1_3_lut_rep_272_4_lut (.A(n8110), .B(select_clk), .C(state_adj_1040[0]), 
         .D(n33447), .Z(n31695)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[17:42])
    defparam i1_3_lut_rep_272_4_lut.init = 16'h0002;
    PFUMX i14614 (.BLUT(n20983), .ALUT(n13), .C0(register_addr[0]), .Z(n6558[6]));
    FD1P3AX reset_count_2573_2574__i1 (.D(n66_adj_1391[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i1.GSR = "ENABLED";
    PFUMX i14611 (.BLUT(n20980), .ALUT(n12), .C0(register_addr[0]), .Z(n20982));
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB encoder_li_pad (.I(encoder_li), .O(encoder_li_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    IB encoder_lb_pad (.I(encoder_lb), .O(encoder_lb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    IB encoder_la_pad (.I(encoder_la), .O(encoder_la_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    IB encoder_ri_pad (.I(encoder_ri), .O(encoder_ri_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    IB encoder_rb_pad (.I(encoder_rb), .O(encoder_rb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    IB encoder_ra_pad (.I(encoder_ra), .O(encoder_ra_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    IB n10608_pad (.I(uart_rx), .O(n10608_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    OB debug_pad_0 (.I(n10608_c), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_1 (.I(n10607), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_6 (.I(n33447), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB motor_pwm_r_pad (.I(GND_net), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    OB expansion5_pad (.I(GND_net), .O(expansion5));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    OB expansion4_pad (.I(GND_net), .O(expansion4));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    OB expansion3_pad (.I(GND_net), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    OB expansion2_pad (.I(GND_net), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion1_pad (.I(GND_net), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    LUT4 i14612_3_lut (.A(Stepper_Y_En_c), .B(div_factor_reg_adj_874[6]), 
         .C(register_addr[1]), .Z(n20983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i14612_3_lut.init = 16'hcaca;
    PFUMX i11332 (.BLUT(n15[3]), .ALUT(n59[3]), .C0(state_adj_1040[1]), 
          .Z(n17735));
    PFUMX i11342 (.BLUT(n15[5]), .ALUT(n59[5]), .C0(state_adj_1040[1]), 
          .Z(n17745));
    PFUMX i11345 (.BLUT(n15[2]), .ALUT(n59[2]), .C0(state_adj_1040[1]), 
          .Z(n17748));
    PFUMX i11350 (.BLUT(n15[4]), .ALUT(n59[4]), .C0(state_adj_1040[1]), 
          .Z(n17753));
    LUT4 i23112_4_lut (.A(reset_count[14]), .B(n29370), .C(reset_count[10]), 
         .D(n29853), .Z(n30)) /* synthesis lut_function=(!(A (B+(C (D))))) */ ;
    defparam i23112_4_lut.init = 16'h5777;
    LUT4 i22706_4_lut (.A(reset_count[9]), .B(n29), .C(n29850), .D(reset_count[6]), 
         .Z(n29853)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i22706_4_lut.init = 16'ha088;
    LUT4 i22704_4_lut (.A(reset_count[5]), .B(n29), .C(n29966), .D(reset_count[4]), 
         .Z(n29850)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i22704_4_lut.init = 16'hfeee;
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB uart_tx_pad (.I(n10607), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    LUT4 i1_4_lut (.A(n33447), .B(state_adj_1182[3]), .C(n24417), .D(state_adj_1182[2]), 
         .Z(n28845)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut.init = 16'h0150;
    LUT4 i1_2_lut (.A(reset_count[9]), .B(reset_count[10]), .Z(n24311)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_adj_478 (.A(reset_count[13]), .B(reset_count[11]), .C(reset_count[12]), 
         .Z(n29370)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_adj_478.init = 16'hfefe;
    LUT4 i2_3_lut_3_lut (.A(n31783), .B(n1294[17]), .C(n1294[20]), .Z(n28025)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i2_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i8_2_lut (.A(state_adj_1040[1]), .B(state_adj_1040[0]), .Z(n7447[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    defparam i8_2_lut.init = 16'h6666;
    LUT4 i23117_4_lut_4_lut (.A(n31783), .B(n4_adj_765), .C(n5613), .D(n1294[14]), 
         .Z(n13568)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i23117_4_lut_4_lut.init = 16'h2a00;
    FD1P3AX reset_count_2573_2574__i2 (.D(n66_adj_1391[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i2.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_479 (.A(register_addr[1]), .B(div_factor_reg_adj_874[9]), 
         .C(steps_reg_adj_875[9]), .D(register_addr[0]), .Z(n99_adj_1262[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_479.init = 16'ha088;
    CCU2D reset_count_2573_2574_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27385), .S0(n66_adj_1391[13]), 
          .S1(n66_adj_1391[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_15.INJECT1_1 = "NO";
    LUT4 i14609_3_lut (.A(control_reg_adj_873[3]), .B(div_factor_reg_adj_874[3]), 
         .C(register_addr[1]), .Z(n20980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i14609_3_lut.init = 16'hcaca;
    FD1P3AX reset_count_2573_2574__i3 (.D(n66_adj_1391[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i4 (.D(n66_adj_1391[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i5 (.D(n66_adj_1391[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i6 (.D(n66_adj_1391[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i7 (.D(n66_adj_1391[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i8 (.D(n66_adj_1391[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i9 (.D(n66_adj_1391[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i10 (.D(n66_adj_1391[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i11 (.D(n66_adj_1391[10]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i12 (.D(n66_adj_1391[11]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i13 (.D(n66_adj_1391[12]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i14 (.D(n66_adj_1391[13]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2573_2574__i15 (.D(n66_adj_1391[14]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574__i15.GSR = "ENABLED";
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.read_value({read_value_adj_956}), 
            .debug_c_c(debug_c_c), .n2669(n2669), .n9093(n9093), .n33450(n33450), 
            .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_957[0]), .n8940(n8940), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .n14252(n14252), .n579(n571_adj_974[0]), .prev_select(prev_select_adj_723), 
            .n31741(n31741), .n33447(n33447), .\register_addr[1] (register_addr[1]), 
            .Stepper_A_M1_c_1(Stepper_A_M1_c_1), .n32(n32_adj_572), .n32_adj_294(n32), 
            .prev_step_clk(prev_step_clk_adj_652), .step_clk(step_clk_adj_651), 
            .n31711(n31711), .n22(n22_adj_571), .n32_adj_295(n32_adj_573), 
            .prev_step_clk_adj_296(prev_step_clk_adj_612), .step_clk_adj_297(step_clk_adj_611), 
            .n31712(n31712), .\register_addr[0] (register_addr[0]), .n22_adj_298(n22), 
            .prev_step_clk_adj_299(prev_step_clk), .n34(n34), .step_clk_adj_300(step_clk), 
            .n31713(n31713), .n24(n24), .n33446(n33446), .n191(n191), 
            .n185(n185), .n33448(n33448), .n33449(n33449), .n33451(n33451), 
            .\read_size[2] (read_size_adj_957[2]), .n29590(n29590), .n31700(n31700), 
            .n33453(n33453), .databus({databus}), .Stepper_A_M2_c_2(Stepper_A_M2_c_2), 
            .Stepper_A_Dir_c(Stepper_A_Dir_c), .Stepper_A_En_c(Stepper_A_En_c), 
            .\control_reg[7] (control_reg_adj_953[7]), .n8885(n8885), .n31784(n31784), 
            .n27905(n27905), .n3700(n3700), .limit_c_3(limit_c_3), .Stepper_A_Step_c(Stepper_A_Step_c), 
            .n8261(n8260[7])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(603[25] 616[45])
    CCU2D reset_count_2573_2574_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27384), .COUT(n27385), .S0(n66_adj_1391[11]), 
          .S1(n66_adj_1391[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2573_2574_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27383), .COUT(n27384), .S0(n66_adj_1391[9]), 
          .S1(n66_adj_1391[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2573_2574_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27382), .COUT(n27383), .S0(n66_adj_1391[7]), 
          .S1(n66_adj_1391[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2573_2574_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27381), .COUT(n27382), .S0(n66_adj_1391[5]), 
          .S1(n66_adj_1391[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_7.INJECT1_1 = "NO";
    GSR GSR_INST (.GSR(VCC_net));
    CCU2D reset_count_2573_2574_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27380), .COUT(n27381), .S0(n66_adj_1391[3]), 
          .S1(n66_adj_1391[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_5.INJECT1_1 = "NO";
    \ClockDividerP_SP(factor=12000000)  encoder_speed_reseter (.GND_net(GND_net), 
            .clk_10Hz(clk_10Hz), .debug_c_c(debug_c_c), .n33448(n33448), 
            .n33447(n33447)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(622[31] 624[67])
    RCPeripheral rc_receiver (.\read_value[18] (read_value_adj_956[18]), .read_value({read_value_adj_996}), 
            .n31719(n31719), .n47(n47_adj_759), .\read_value[18]_adj_91 (read_value_adj_864[18]), 
            .n6(n6_adj_802), .n31703(n31703), .databus_out({databus_out}), 
            .rw(rw), .\read_value[18]_adj_92 (read_value_adj_916[18]), .read_value_adj_293({read_value}), 
            .n31716(n31716), .n46(n46), .n3(n3_adj_809), .databus({databus}), 
            .\read_value[17]_adj_125 (read_value_adj_956[17]), .\read_value[17]_adj_126 (read_value_adj_864[17]), 
            .n6_adj_127(n6_adj_810), .\read_value[6]_adj_128 (read_value_adj_876[6]), 
            .n31733(n31733), .n33446(n33446), .\read_value[17]_adj_129 (read_value_adj_916[17]), 
            .\read_value[6]_adj_130 (read_value_adj_864[6]), .n3_adj_131(n3_adj_807), 
            .\select[7] (select[7]), .\read_value[16]_adj_132 (read_value_adj_956[16]), 
            .\read_value[16]_adj_133 (read_value_adj_864[16]), .n6_adj_134(n6_adj_808), 
            .\read_value[16]_adj_135 (read_value_adj_916[16]), .n3_adj_136(n3_adj_798), 
            .\read_value[15]_adj_137 (read_value_adj_956[15]), .\read_value[15]_adj_138 (read_value_adj_864[15]), 
            .n6_adj_139(n6_adj_724), .\read_value[15]_adj_140 (read_value_adj_916[15]), 
            .\register_addr[0] (register_addr[0]), .n8(n8_adj_784), .\read_value[7]_adj_141 (read_value_adj_876[7]), 
            .n3_adj_142(n3_adj_796), .\read_value[14]_adj_143 (read_value_adj_956[14]), 
            .\read_value[14]_adj_144 (read_value_adj_864[14]), .n6_adj_145(n6_adj_797), 
            .n8_adj_146(n8), .\read_value[14]_adj_147 (read_value_adj_916[14]), 
            .n3_adj_148(n3_adj_789), .\read_value[13]_adj_149 (read_value_adj_956[13]), 
            .\read_value[13]_adj_150 (read_value_adj_864[13]), .n6_adj_151(n6_adj_791), 
            .\read_value[13]_adj_152 (read_value_adj_916[13]), .\read_value[7]_adj_153 (read_value_adj_864[7]), 
            .n3_adj_154(n3_adj_786), .n3_adj_155(n3_adj_768), .\read_value[31]_adj_156 (read_value_adj_956[31]), 
            .\read_value[12]_adj_157 (read_value_adj_956[12]), .\read_value[12]_adj_158 (read_value_adj_864[12]), 
            .n6_adj_159(n6_adj_788), .\read_value[31]_adj_160 (read_value_adj_864[31]), 
            .n6_adj_161(n6_adj_767), .\read_value[12]_adj_162 (read_value_adj_916[12]), 
            .\read_value[31]_adj_163 (read_value_adj_916[31]), .n3_adj_164(n3_adj_790), 
            .\read_value[11]_adj_165 (read_value_adj_956[11]), .\read_value[11]_adj_166 (read_value_adj_864[11]), 
            .n6_adj_167(n6_adj_792), .\read_value[11]_adj_168 (read_value_adj_916[11]), 
            .\register_addr[2] (register_addr[2]), .\register_addr[1] (register_addr[1]), 
            .n3_adj_169(n3_adj_785), .\read_value[10]_adj_170 (read_value_adj_956[10]), 
            .\read_value[10]_adj_171 (read_value_adj_864[10]), .n6_adj_172(n6_adj_787), 
            .n3_adj_173(n3_adj_778), .\read_value[30]_adj_174 (read_value_adj_956[30]), 
            .\read_value[30]_adj_175 (read_value_adj_864[30]), .n6_adj_176(n6_adj_775), 
            .\read_value[10]_adj_177 (read_value_adj_916[10]), .\read_value[30]_adj_178 (read_value_adj_916[30]), 
            .n3_adj_179(n3_adj_831), .\read_value[29]_adj_180 (read_value_adj_956[29]), 
            .\read_value[29]_adj_181 (read_value_adj_864[29]), .n6_adj_182(n6_adj_824), 
            .\read_value[29]_adj_183 (read_value_adj_916[29]), .n3_adj_184(n3_adj_794), 
            .\read_value[9]_adj_185 (read_value_adj_956[9]), .n3_adj_186(n3_adj_648), 
            .\read_value[28]_adj_187 (read_value_adj_956[28]), .\read_value[9]_adj_188 (read_value_adj_864[9]), 
            .n6_adj_189(n6_adj_795), .\read_value[28]_adj_190 (read_value_adj_864[28]), 
            .n6_adj_191(n6), .\read_value[28]_adj_192 (read_value_adj_916[28]), 
            .\read_value[9]_adj_193 (read_value_adj_916[9]), .n3_adj_194(n3_adj_817), 
            .\read_value[27]_adj_195 (read_value_adj_956[27]), .n3_adj_196(n3), 
            .\read_value[27]_adj_197 (read_value_adj_864[27]), .n6_adj_198(n6_adj_818), 
            .\read_value[27]_adj_199 (read_value_adj_916[27]), .\read_value[8]_adj_200 (read_value_adj_956[8]), 
            .\read_value[8]_adj_201 (read_value_adj_864[8]), .n6_adj_202(n6_adj_793), 
            .\read_value[8]_adj_203 (read_value_adj_916[8]), .n3_adj_204(n3_adj_822), 
            .\read_value[26]_adj_205 (read_value_adj_956[26]), .\read_value[26]_adj_206 (read_value_adj_864[26]), 
            .n6_adj_207(n6_adj_816), .\read_value[26]_adj_208 (read_value_adj_916[26]), 
            .n3_adj_209(n3_adj_820), .\read_value[25]_adj_210 (read_value_adj_956[25]), 
            .\read_value[25]_adj_211 (read_value_adj_864[25]), .n6_adj_212(n6_adj_821), 
            .\read_value[25]_adj_213 (read_value_adj_916[25]), .\read_size[0] (read_size_adj_858[0]), 
            .\read_size[0]_adj_214 (read_size_adj_1006[0]), .\select[2] (select[2]), 
            .n31780(n31780), .n9(n9_adj_766), .n29694(n29694), .n14(n14), 
            .n3_adj_215(n3_adj_815), .\select[4] (select[4]), .\read_size[0]_adj_216 (read_size_adj_997[0]), 
            .n55(n55), .n31762(n31762), .n10(n10), .read_size({read_size}), 
            .n31732(n31732), .\select[1] (select[1]), .\read_size[0]_adj_218 (read_size_adj_917[0]), 
            .n31741(n31741), .n6_adj_219(n6_adj_829), .\read_size[2]_adj_220 (read_size_adj_957[2]), 
            .\reg_size[2] (reg_size[2]), .n9_adj_221(n9_adj_825), .\read_size[2]_adj_222 (read_size_adj_917[2]), 
            .\read_value[24]_adj_223 (read_value_adj_956[24]), .\read_value[24]_adj_224 (read_value_adj_864[24]), 
            .n6_adj_225(n6_adj_819), .\read_size[2]_adj_226 (read_size_adj_1006[2]), 
            .n2(n2_adj_773), .\read_value[5]_adj_227 (read_value_adj_956[5]), 
            .n5(n5_adj_774), .n8_adj_228(n8_adj_772), .\read_value[24]_adj_229 (read_value_adj_916[24]), 
            .n3_adj_230(n3_adj_813), .\read_value[23]_adj_231 (read_value_adj_956[23]), 
            .\read_value[23]_adj_232 (read_value_adj_864[23]), .n6_adj_233(n6_adj_814), 
            .n2_adj_234(n2_adj_779), .\read_value[23]_adj_235 (read_value_adj_916[23]), 
            .\read_value[5]_adj_236 (read_value_adj_876[5]), .\read_value[6]_adj_237 (read_value_adj_956[6]), 
            .n5_adj_238(n5_adj_780), .n3_adj_239(n3_adj_811), .\read_value[5]_adj_240 (read_value_adj_864[5]), 
            .\read_value[22]_adj_241 (read_value_adj_956[22]), .\read_value[22]_adj_242 (read_value_adj_864[22]), 
            .n6_adj_243(n6_adj_812), .\read_value[22]_adj_244 (read_value_adj_916[22]), 
            .n3_adj_245(n3_adj_803), .\read_value[21]_adj_246 (read_value_adj_956[21]), 
            .\read_value[21]_adj_247 (read_value_adj_864[21]), .n6_adj_248(n6_adj_804), 
            .\read_value[21]_adj_249 (read_value_adj_916[21]), .n3_adj_250(n3_adj_799), 
            .n31841(n31841), .\sendcount[1] (sendcount[1]), .n12795(n12795), 
            .\read_value[20]_adj_251 (read_value_adj_956[20]), .\read_value[20]_adj_252 (read_value_adj_864[20]), 
            .n6_adj_253(n6_adj_801), .\read_value[20]_adj_254 (read_value_adj_916[20]), 
            .n2_adj_255(n2_adj_776), .n3_adj_256(n3_adj_805), .\read_value[19]_adj_257 (read_value_adj_956[19]), 
            .\read_value[19]_adj_258 (read_value_adj_864[19]), .n6_adj_259(n6_adj_806), 
            .\read_value[4]_adj_260 (read_value_adj_956[4]), .n5_adj_261(n5_adj_649), 
            .n8_adj_262(n8_adj_781), .\read_value[19]_adj_263 (read_value_adj_916[19]), 
            .n3_adj_264(n3_adj_800), .n8_adj_265(n8_adj_777), .\read_value[4]_adj_266 (read_value_adj_876[4]), 
            .\read_value[4]_adj_267 (read_value_adj_864[4]), .n2_adj_268(n2_adj_769), 
            .\read_value[3]_adj_269 (read_value_adj_956[3]), .n5_adj_270(n5_adj_770), 
            .n8_adj_271(n8_adj_771), .\read_value[3]_adj_272 (read_value_adj_876[3]), 
            .\read_value[3]_adj_273 (read_value_adj_864[3]), .\read_value[7]_adj_274 (read_value_adj_956[7]), 
            .n5_adj_275(n5_adj_783), .n29738(n29738), .n2_adj_276(n2), 
            .\read_value[2]_adj_277 (read_value_adj_956[2]), .n5_adj_278(n5_adj_570), 
            .n8_adj_279(n8_adj_823), .\read_value[2]_adj_280 (read_value_adj_876[2]), 
            .\read_value[2]_adj_281 (read_value_adj_864[2]), .n1(n1), .n5_adj_282(n5), 
            .\read_value[0]_adj_283 (read_value_adj_864[0]), .n2_adj_284(n2_adj_763), 
            .\read_value[0]_adj_285 (read_value_adj_876[0]), .\read_value[1]_adj_286 (read_value_adj_876[1]), 
            .n4(n4), .n2_adj_287(n2_adj_782), .\read_value[1]_adj_288 (read_value_adj_1005[1]), 
            .n31746(n31746), .n2_adj_289(n2_adj_827), .\read_value[0]_adj_290 (read_value_adj_956[0]), 
            .n5_adj_291(n5_adj_826), .GND_net(GND_net), .debug_c_c(debug_c_c), 
            .n31694(n31694), .rc_ch8_c(rc_ch8_c), .n27918(n27918), .n30160(n30160), 
            .n30216(n30216), .n13719(n13719), .rc_ch7_c(rc_ch7_c), .n27933(n27933), 
            .n30195(n30195), .n14176(n14176), .n30205(n30205), .rc_ch4_c(rc_ch4_c), 
            .n27937(n27937), .n30182(n30182), .n14182(n14182), .n30191(n30191), 
            .n30197(n30197), .rc_ch3_c(rc_ch3_c), .n27924(n27924), .n14183(n14183), 
            .n30189(n30189), .n30186(n30186), .rc_ch2_c(rc_ch2_c), .n27915(n27915), 
            .n14186(n14186), .n30218(n30218), .n29930(n29930), .n14187(n14187), 
            .n9_adj_292(n9), .rc_ch1_c(rc_ch1_c), .n30152(n30152), .n30184(n30184), 
            .n27912(n27912)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(670[15] 682[41])
    CCU2D reset_count_2573_2574_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27379), .COUT(n27380), .S0(n66_adj_1391[1]), 
          .S1(n66_adj_1391[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2573_2574_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2573_2574_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27379), .S1(n66_adj_1391[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2573_2574_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2573_2574_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2573_2574_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2573_2574_add_4_1.INJECT1_1 = "NO";
    \ProtocolInterface(baud_div=12)  protocol_interface (.debug_c_c(debug_c_c), 
            .n33455(n33455), .\select[7] (select[7]), .\select[1] (select[1]), 
            .\select[4] (select[4]), .\select[2] (select[2]), .databus_out({databus_out}), 
            .n13568(n13568), .\read_value[6] (read_value_adj_916[6]), .n33446(n33446), 
            .n2(n2_adj_779), .register_addr({Open_31, Open_32, register_addr[5], 
            Open_33, Open_34, register_addr[2], Open_35, register_addr[0]}), 
            .n31751(n31751), .\read_value[3] (read_value_adj_916[3]), .rw(rw), 
            .n2_adj_43(n2_adj_769), .\register[2][0] (\register[2] [0]), 
            .\register_addr[3] (register_addr[3]), .n31716(n31716), .\register_addr[1] (register_addr[1]), 
            .\steps_reg[5] (steps_reg_adj_875[5]), .n14(n14_adj_830), .\read_value[4] (read_value_adj_916[4]), 
            .n2_adj_44(n2_adj_776), .n31827(n31827), .n27707(n27707), 
            .n31720(n31720), .n33447(n33447), .n14124(n14124), .\read_value[7] (read_value_adj_916[7]), 
            .n2_adj_45(n2_adj_782), .n1306(n1294[20]), .\read_value[2] (read_value_adj_916[2]), 
            .n2_adj_46(n2), .n1309(n1294[17]), .n1312(n1294[14]), .\read_value[1] (read_value_adj_916[1]), 
            .n2_adj_47(n2_adj_763), .\read_value[0] (read_value_adj_916[0]), 
            .n2_adj_48(n2_adj_827), .\read_value[5] (read_value_adj_916[5]), 
            .n2_adj_49(n2_adj_773), .n31717(n31717), .n31867(n31867), 
            .n31698(n31698), .n191(n191), .n29590(n29590), .n31699(n31699), 
            .n13671(n13671), .n31705(n31705), .n8940(n8940), .\sendcount[1] (sendcount[1]), 
            .prev_select(prev_select_adj_687), .n2658(n2658), .n21(n21), 
            .n29452(n29452), .n185(n185), .n14252(n14252), .\register_addr[4] (register_addr[4]), 
            .n31746(n31746), .debug_c_7(debug_c_7), .n13757(n13757), .n31779(n31779), 
            .n29552(n29552), .n47(n47_adj_759), .\read_size[2] (read_size_adj_997[2]), 
            .n6(n6_adj_829), .n31739(n31739), .\read_value[1]_adj_50 (read_value_adj_864[1]), 
            .n4(n4), .n3970(n3970), .n78(n78_adj_832), .n31763(n31763), 
            .\read_value[19] (read_value_adj_876[19]), .n3(n3_adj_805), 
            .\read_value[20] (read_value_adj_876[20]), .n3_adj_51(n3_adj_799), 
            .\read_size[2]_adj_52 (read_size_adj_877[2]), .n31832(n31832), 
            .\read_value[21] (read_value_adj_876[21]), .n3_adj_53(n3_adj_803), 
            .prev_select_adj_54(prev_select_adj_609), .n14172(n14172), .\read_value[22] (read_value_adj_876[22]), 
            .n3_adj_55(n3_adj_811), .\read_value[23] (read_value_adj_876[23]), 
            .n3_adj_56(n3_adj_813), .\read_value[24] (read_value_adj_876[24]), 
            .n3_adj_57(n3_adj_815), .\read_value[25] (read_value_adj_876[25]), 
            .n3_adj_58(n3_adj_820), .\read_value[26] (read_value_adj_876[26]), 
            .n3_adj_59(n3_adj_822), .\read_value[27] (read_value_adj_876[27]), 
            .n3_adj_60(n3_adj_817), .\read_value[28] (read_value_adj_876[28]), 
            .n3_adj_61(n3_adj_648), .\read_value[29] (read_value_adj_876[29]), 
            .n3_adj_62(n3_adj_831), .\read_value[30] (read_value_adj_876[30]), 
            .n3_adj_63(n3_adj_778), .n31741(n31741), .\read_value[31] (read_value_adj_876[31]), 
            .n3_adj_64(n3_adj_768), .\read_value[18] (read_value_adj_876[18]), 
            .n3_adj_65(n3_adj_800), .\read_value[17] (read_value_adj_876[17]), 
            .n3_adj_66(n3_adj_809), .\read_value[16] (read_value_adj_876[16]), 
            .n3_adj_67(n3_adj_807), .\read_value[15] (read_value_adj_876[15]), 
            .n3_adj_68(n3_adj_798), .\read_value[14] (read_value_adj_876[14]), 
            .n3_adj_69(n3_adj_796), .\read_value[13] (read_value_adj_876[13]), 
            .n3_adj_70(n3_adj_789), .n31783(n31783), .databus({databus}), 
            .\read_value[12] (read_value_adj_876[12]), .n3_adj_71(n3_adj_786), 
            .\read_value[11] (read_value_adj_876[11]), .n3_adj_72(n3_adj_790), 
            .\read_value[10] (read_value_adj_876[10]), .n3_adj_73(n3_adj_785), 
            .n28025(n28025), .n33445(n33445), .n33457(n33457), .n28937(n28937), 
            .n31780(n31780), .\read_value[9] (read_value_adj_876[9]), .n3_adj_74(n3_adj_794), 
            .n22093(n22093), .\read_value[8] (read_value_adj_876[8]), .n3_adj_75(n3), 
            .n31762(n31762), .prev_select_adj_76(prev_select), .n29823(n29823), 
            .n31703(n31703), .n31718(n31718), .n31774(n31774), .n14022(n14022), 
            .n16046(n16046), .n16045(n16045), .n24748(n24748), .n250(n249[2]), 
            .\read_value[1]_adj_77 (read_value_adj_956[1]), .n1(n1), .n29738(n29738), 
            .\steps_reg[6] (steps_reg_adj_875[6]), .n13(n13), .n31724(n31724), 
            .n12795(n12795), .n9(n9_adj_766), .n14_adj_78(n14), .n10(n10), 
            .\reg_size[2] (reg_size[2]), .n31841(n31841), .n106(n106), 
            .\control_reg[7] (control_reg_adj_873[7]), .n8243(n8242[7]), 
            .\read_size[0] (read_size_adj_957[0]), .\read_size[0]_adj_79 (read_size_adj_865[0]), 
            .n55(n55), .\read_size[2]_adj_80 (read_size_adj_865[2]), .n9_adj_81(n9_adj_825), 
            .\control_reg[7]_adj_82 (control_reg[7]), .n1_adj_83(n1_adj_764), 
            .n5613(n5613), .n31722(n31722), .n13779(n13779), .n31707(n31707), 
            .n31785(n31785), .n14084(n14084), .\read_size[0]_adj_84 (read_size_adj_877[0]), 
            .n29694(n29694), .n13476(n13476), .\control_reg[7]_adj_85 (control_reg_adj_913[7]), 
            .n8252(n8251[7]), .n4_adj_86(n4_adj_765), .\control_reg[7]_adj_87 (control_reg_adj_953[7]), 
            .n8261(n8260[7]), .n31733(n31733), .\steps_reg[3] (steps_reg_adj_875[3]), 
            .n12(n12), .\arm_select[0] (arm_select[0]), .n31727(n31727), 
            .prev_select_adj_88(prev_select_adj_647), .n3883(n3883), .n9089(n9089), 
            .n24720(n24720), .n24690(n24690), .n13606(n13606), .n89(n89_adj_833), 
            .n31732(n31732), .n3786(n3786), .n31700(n31700), .n3700(n3700), 
            .n8885(n8885), .debug_c_2(debug_c_2), .debug_c_3(debug_c_3), 
            .debug_c_4(debug_c_4), .debug_c_5(debug_c_5), .n31701(n31701), 
            .n24729(n24729), .n31708(n31708), .prev_select_adj_89(prev_select_adj_723), 
            .n31715(n31715), .n31719(n31719), .n10607(n10607), .GND_net(GND_net), 
            .n10608_c(n10608_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[26] 485[57])
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.read_value({read_value_adj_916}), 
            .debug_c_c(debug_c_c), .n2658(n2658), .VCC_net(VCC_net), .GND_net(GND_net), 
            .Stepper_Z_nFault_c(Stepper_Z_nFault_c), .n33450(n33450), .\read_size[0] (read_size_adj_917[0]), 
            .n24720(n24720), .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n13779(n13779), 
            .n579(n571_adj_974[0]), .prev_step_clk(prev_step_clk_adj_652), 
            .step_clk(step_clk_adj_651), .n13757(n13757), .prev_select(prev_select_adj_687), 
            .n31732(n31732), .n31707(n31707), .n33448(n33448), .databus({databus}), 
            .n33449(n33449), .\control_reg[7] (control_reg_adj_913[7]), 
            .n31722(n31722), .Stepper_Z_En_c(Stepper_Z_En_c), .Stepper_Z_Dir_c(Stepper_Z_Dir_c), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), 
            .n27902(n27902), .n9089(n9089), .\register_addr[0] (register_addr[0]), 
            .n32(n32), .n22(n22_adj_571), .n31711(n31711), .\register_addr[1] (register_addr[1]), 
            .\read_size[2] (read_size_adj_917[2]), .n24690(n24690), .n33451(n33451), 
            .n33452(n33452), .n3786(n3786), .limit_c_2(limit_c_2), .n33447(n33447), 
            .Stepper_Z_Step_c(Stepper_Z_Step_c), .n8252(n8251[7])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(588[25] 601[45])
    VLO i1 (.Z(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i1_3_lut (.A(n33447), .B(limit_latched), .C(prev_limit_latched), 
         .Z(n10675)) /* synthesis lut_function=(A+!((C)+!B)) */ ;
    defparam i1_3_lut.init = 16'haeae;
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.\read_size[2] (read_size_adj_865[2]), 
            .debug_c_c(debug_c_c), .n13671(n13671), .n31720(n31720), .GND_net(GND_net), 
            .n33451(n33451), .databus({databus}), .n3970(n3970), .n33450(n33450), 
            .step_clk(step_clk), .n34(n34), .prev_step_clk(prev_step_clk), 
            .\read_size[0] (read_size_adj_865[0]), .n106(n106), .Stepper_X_M0_c_0(Stepper_X_M0_c_0), 
            .n14172(n14172), .n579(n571_adj_974[0]), .limit_latched(limit_latched), 
            .prev_limit_latched(prev_limit_latched), .n14124(n14124), .prev_select(prev_select_adj_609), 
            .\arm_select[0] (arm_select[0]), .n29552(n29552), .\register_addr[0] (register_addr[0]), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\register_addr[1] (register_addr[1]), 
            .n24(n24), .n31713(n31713), .n31702(n31702), .n33453(n33453), 
            .n608(n580[4]), .n610(n580[2]), .\control_reg[7] (control_reg[7]), 
            .n31701(n31701), .n10675(n10675), .Stepper_X_En_c(Stepper_X_En_c), 
            .Stepper_X_Dir_c(Stepper_X_Dir_c), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), 
            .n27910(n27910), .VCC_net(VCC_net), .Stepper_X_nFault_c(Stepper_X_nFault_c), 
            .read_value({read_value_adj_864}), .n31705(n31705), .limit_c_0(limit_c_0), 
            .n1(n1_adj_764), .Stepper_X_Step_c(Stepper_X_Step_c), .n33447(n33447), 
            .n33448(n33448)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(558[25] 571[45])
    LUT4 i23074_2_lut (.A(int_step), .B(control_reg_adj_873[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i23074_2_lut.init = 16'h9999;
    LUT4 m1_lut (.Z(n33445)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    LUT4 i3_4_lut (.A(n31818), .B(n31797), .C(n31798), .D(n9848), .Z(n27884)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i3_4_lut.init = 16'h1000;
    ClockDivider_U10 pwm_clk_div (.n33447(n33447), .n7485(n7485), .n30160(n30160), 
            .n13719(n13719), .debug_c_c(debug_c_c), .n241(n241), .n30205(n30205), 
            .n14176(n14176), .n30191(n30191), .n14182(n14182), .n30189(n30189), 
            .n14183(n14183), .n30186(n30186), .n14186(n14186), .n29930(n29930), 
            .n9(n9), .n30184(n30184), .n14187(n14187), .n30182(n30182), 
            .n27937(n27937), .n30195(n30195), .n27933(n27933), .n30197(n30197), 
            .n27924(n27924), .n30216(n30216), .n27918(n27918), .n31694(n31694), 
            .n30218(n30218), .n27915(n27915), .n30152(n30152), .n27912(n27912), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(518[15] 521[41])
    EncoderPeripheral_U11 left_encoder (.\read_size[0] (read_size_adj_997[0]), 
            .n31762(n31762), .n24748(n24748), .read_value({read_value_adj_996}), 
            .n33457(n33457), .n31717(n31717), .encoder_la_c(encoder_la_c), 
            .\register_addr[0] (register_addr[0]), .encoder_lb_c(encoder_lb_c), 
            .\read_size[2] (read_size_adj_997[2]), .n250(n249[2]), .encoder_li_c(encoder_li_c), 
            .n33447(n33447), .clk_10Hz(clk_10Hz), .n31759(n31759), .n4144(n4137[25]), 
            .n47(n99_adj_1259[25]), .debug_c_c(debug_c_c), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(646[20] 656[47])
    EncoderPeripheral right_encoder (.n31780(n31780), .n33457(n33457), .\read_size[0] (read_size_adj_1006[0]), 
            .n24748(n24748), .encoder_ri_c(encoder_ri_c), .\register_addr[0] (register_addr[0]), 
            .encoder_rb_c(encoder_rb_c), .encoder_ra_c(encoder_ra_c), .rw(rw), 
            .n6(n6_adj_821), .n6_adj_14(n6_adj_806), .n6_adj_15(n6_adj_819), 
            .n6_adj_16(n6_adj_814), .n6_adj_17(n6_adj_812), .n6_adj_18(n6_adj_804), 
            .n6_adj_19(n6_adj_801), .n6_adj_20(n6_adj_802), .n6_adj_21(n6_adj_810), 
            .n6_adj_22(n6_adj_808), .n6_adj_23(n6_adj_724), .n6_adj_24(n6_adj_797), 
            .n6_adj_25(n6_adj_791), .n6_adj_26(n6_adj_788), .n6_adj_27(n6_adj_792), 
            .n6_adj_28(n6_adj_787), .n6_adj_29(n6_adj_795), .n6_adj_30(n6_adj_793), 
            .\read_value[1] (read_value_adj_1005[1]), .n31717(n31717), .n31708(n31708), 
            .\read_size[2] (read_size_adj_1006[2]), .n250(n249[2]), .n8(n8_adj_823), 
            .n8_adj_31(n8), .n6_adj_32(n6_adj_767), .n6_adj_33(n6_adj_775), 
            .n6_adj_34(n6_adj_824), .n6_adj_35(n6), .n6_adj_36(n6_adj_818), 
            .n6_adj_37(n6_adj_816), .n8_adj_38(n8_adj_784), .n8_adj_39(n8_adj_781), 
            .n8_adj_40(n8_adj_772), .n8_adj_41(n8_adj_777), .n8_adj_42(n8_adj_771), 
            .debug_c_c(debug_c_c), .n31759(n31759), .n47(n99_adj_1259[25]), 
            .GND_net(GND_net), .n4144(n4137[25]), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(657[20] 667[47])
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .VCC_net(VCC_net), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .n33450(n33450), .\read_size[0] (read_size_adj_877[0]), .n14194(n14194), 
            .n78(n78_adj_832), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), .n89(n89_adj_833), 
            .n579(n571_adj_974[0]), .prev_step_clk(prev_step_clk_adj_612), 
            .step_clk(step_clk_adj_611), .n14084(n14084), .prev_select(prev_select_adj_647), 
            .n31727(n31727), .\steps_reg[9] (steps_reg_adj_875[9]), .\steps_reg[5] (steps_reg_adj_875[5]), 
            .\steps_reg[6] (steps_reg_adj_875[6]), .\steps_reg[3] (steps_reg_adj_875[3]), 
            .n32(n32_adj_573), .\register_addr[0] (register_addr[0]), .n27893(n27893), 
            .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), .int_step(int_step), .n22(n22), 
            .n31712(n31712), .n31724(n31724), .n33448(n33448), .databus({databus}), 
            .n33451(n33451), .n33452(n33452), .\div_factor_reg[9] (div_factor_reg_adj_874[9]), 
            .\div_factor_reg[6] (div_factor_reg_adj_874[6]), .\div_factor_reg[5] (div_factor_reg_adj_874[5]), 
            .\div_factor_reg[3] (div_factor_reg_adj_874[3]), .\control_reg[7] (control_reg_adj_873[7]), 
            .n13606(n13606), .Stepper_Y_En_c(Stepper_Y_En_c), .Stepper_Y_Dir_c(Stepper_Y_Dir_c), 
            .\control_reg[3] (control_reg_adj_873[3]), .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), 
            .\read_size[2] (read_size_adj_877[2]), .n33453(n33453), .read_value({read_value_adj_876}), 
            .\register_addr[1] (register_addr[1]), .n8243(n8242[7]), .n3883(n3883), 
            .n33447(n33447), .limit_c_1(limit_c_1), .n31785(n31785), .\register_addr[3] (register_addr[3]), 
            .\register_addr[2] (register_addr[2]), .n79(n99_adj_1262[9]), 
            .n6584(n6558[6]), .n20993(n20993), .n20982(n20982)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(573[25] 586[45])
    SabertoothSerialPeripheral motor_serial (.debug_c_c(debug_c_c), .n13476(n13476), 
            .n31699(n31699), .n33451(n33451), .\databus[6] (databus[6]), 
            .\databus[5] (databus[5]), .\databus[4] (databus[4]), .\databus[3] (databus[3]), 
            .\databus[2] (databus[2]), .\register[1][1] (\register[1]_adj_855 [1]), 
            .\databus[1] (databus[1]), .\databus[0] (databus[0]), .\register[0] ({\register[0]_adj_856 [7], 
            Open_36, Open_37, Open_38, Open_39, Open_40, Open_41, 
            Open_42}), .n22093(n22093), .n31698(n31698), .\register[0][1] (\register[0]_adj_856 [1]), 
            .\read_size[0] (read_size_adj_858[0]), .n106(n106), .n33450(n33450), 
            .\select[2] (select[2]), .n31867(n31867), .n33447(n33447), 
            .\register_addr[0] (register_addr[0]), .n31832(n31832), .n21959(n21959), 
            .n31796(n31796), .n21892(n21892), .n31818(n31818), .rw(rw), 
            .n5(n5_adj_826), .n5_adj_5(n5), .n5_adj_6(n5_adj_570), .n5_adj_7(n5_adj_770), 
            .n5_adj_8(n5_adj_649), .n5_adj_9(n5_adj_774), .n5_adj_10(n5_adj_780), 
            .n5_adj_11(n5_adj_783), .\state[0] (state_adj_1040[0]), .n17748(n17748), 
            .n17735(n17735), .n17753(n17753), .n17745(n17745), .GND_net(GND_net), 
            .n31695(n31695), .\state[1] (state_adj_1040[1]), .n27884(n27884), 
            .n31(n31), .n21729(n21729), .n31797(n31797), .n19(n19), 
            .n9848(n9848), .n7450(n7447[1]), .n44(n15[3]), .n88(n59[3]), 
            .n42(n15[5]), .n86(n59[5]), .n45(n15[2]), .n89(n59[2]), 
            .n43(n15[4]), .n87(n59[4]), .\state[2] (state_adj_1182[2]), 
            .n8110(n8110), .select_clk(select_clk), .\reset_count[14] (reset_count[14]), 
            .\reset_count[12] (reset_count[12]), .\reset_count[13] (reset_count[13]), 
            .n31783(n31783), .n31751(n31751), .n24311(n24311), .n29370(n29370), 
            .n31784(n31784), .\state[3] (state_adj_1182[3]), .n24417(n24417), 
            .n33449(n33449), .n33453(n33453), .n33455(n33455), .n31237(n31237), 
            .\reset_count[0] (reset_count[0]), .\reset_count[3] (reset_count[3]), 
            .\reset_count[2] (reset_count[2]), .\reset_count[1] (reset_count[1]), 
            .n29966(n29966), .n7485(n7485), .n241(n241), .n29(n29), 
            .\reset_count[5] (reset_count[5]), .\reset_count[6] (reset_count[6]), 
            .\reset_count[4] (reset_count[4]), .\reset_count[11] (reset_count[11]), 
            .\reset_count[8] (reset_count[8]), .\reset_count[7] (reset_count[7]), 
            .n14424(n14424), .n33448(n33448), .\databus[7] (databus[7]), 
            .n31779(n31779), .n191(n191), .n31715(n31715), .n9093(n9093), 
            .prev_select(prev_select_adj_723), .n31774(n31774), .\select[4] (select[4]), 
            .n2669(n2669), .n28845(n28845), .n33452(n33452), .n31739(n31739), 
            .\register_addr[1] (register_addr[1]), .n610(n580[2]), .n608(n580[4]), 
            .\register_addr[4] (register_addr[4]), .prev_select_adj_12(prev_select_adj_609), 
            .n31763(n31763), .n13671(n13671), .prev_select_adj_13(prev_select_adj_647), 
            .n14194(n14194), .n579(n571_adj_974[0]), .motor_pwm_l_c(motor_pwm_l_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(508[29] 516[56])
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (\register[2] , debug_c_c, n33450, read_size, 
            n14022, n24748, prev_select, \select[1] , n33449, n33446, 
            n46, read_value, n28937, GND_net, n33448, \databus[1] , 
            \register_addr[1] , n31739, \register_addr[0] , n27707, 
            n31827, n31702, rw, n33447, n29823, n24729, n31720, 
            n31832, \control_reg[7] , n27893, n32, \control_reg[7]_adj_301 , 
            n27905, n32_adj_302, n21959, \register[1][1] , n31796, 
            signal_light_c, \control_reg[7]_adj_303 , n27902, n32_adj_304, 
            \control_reg[7]_adj_305 , n27910, n34, n21892, \register[0][1] , 
            n31797, \register[0][7] , n31798, n21729, n31, \state[0] , 
            n19, \register_addr[2] , n29738, n21, n31779, \register_addr[5] , 
            \register_addr[4] , xbee_pause_c, n16046, n16045, n31718, 
            n29452) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[2] ;
    input debug_c_c;
    input n33450;
    output [2:0]read_size;
    output n14022;
    input n24748;
    output prev_select;
    input \select[1] ;
    input n33449;
    input n33446;
    output n46;
    output [31:0]read_value;
    input n28937;
    input GND_net;
    input n33448;
    input \databus[1] ;
    input \register_addr[1] ;
    input n31739;
    input \register_addr[0] ;
    input n27707;
    input n31827;
    output n31702;
    input rw;
    input n33447;
    input n29823;
    input n24729;
    input n31720;
    output n31832;
    input \control_reg[7] ;
    input n27893;
    output n32;
    input \control_reg[7]_adj_301 ;
    input n27905;
    output n32_adj_302;
    input n21959;
    input \register[1][1] ;
    output n31796;
    output signal_light_c;
    input \control_reg[7]_adj_303 ;
    input n27902;
    output n32_adj_304;
    input \control_reg[7]_adj_305 ;
    input n27910;
    output n34;
    input n21892;
    input \register[0][1] ;
    output n31797;
    input \register[0][7] ;
    output n31798;
    output n21729;
    input n31;
    input \state[0] ;
    output n19;
    input \register_addr[2] ;
    input n29738;
    output n21;
    input n31779;
    input \register_addr[5] ;
    input \register_addr[4] ;
    input xbee_pause_c;
    input n16046;
    input n16045;
    input n31718;
    input n29452;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n31831;
    wire [31:0]n100;
    
    wire prev_clk_1Hz, clk_1Hz;
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n178;
    wire [31:0]\register[2]_c ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n9030, n9075, n27226, n27225, n27224, n27223, n27222, 
        n27221, force_pause, n28621, n27220, n27219, n27218, n29504, 
        n27217, n27216, n27215, n27214, n27213, n29503, n27212, 
        n27211, n29506, n29501, n29505, n29499, n29500, n29497, 
        n29486, n29509, n29496, n29491, n29489, n29487, n29507, 
        n28853, n29495, n29510, n29494, n29508, n29490, n29493, 
        n29484, n29483, n29502, n29488, n29485, n29492, n29498, 
        n29739, n24, n28729;
    
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n31831), .CD(n33450), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n24748), .SP(n14022), .CK(debug_c_c), 
            .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_149 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_clk_1Hz_149.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_150 (.D(n178), .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam xbee_pause_latched_150.GSR = "ENABLED";
    FD1S3AX prev_select_148 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_select_148.GSR = "ENABLED";
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n9030), .CD(n33449), 
            .CK(debug_c_c), .Q(\register[2]_c [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n9030), .CD(n33449), .CK(debug_c_c), 
            .Q(\register[2]_c [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n9030), .CD(n33450), .CK(debug_c_c), 
            .Q(\register[2]_c [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    LUT4 i14_2_lut (.A(\select[1] ), .B(n33446), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam i14_2_lut.init = 16'h8888;
    FD1P3IX read_value__i0 (.D(n28937), .SP(n14022), .CD(n9075), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i0.GSR = "ENABLED";
    CCU2D add_134_33 (.A0(\register[2]_c [31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27226), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_33.INIT0 = 16'h5aaa;
    defparam add_134_33.INIT1 = 16'h0000;
    defparam add_134_33.INJECT1_0 = "NO";
    defparam add_134_33.INJECT1_1 = "NO";
    CCU2D add_134_31 (.A0(\register[2]_c [29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27225), .COUT(n27226), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_31.INIT0 = 16'h5aaa;
    defparam add_134_31.INIT1 = 16'h5aaa;
    defparam add_134_31.INJECT1_0 = "NO";
    defparam add_134_31.INJECT1_1 = "NO";
    CCU2D add_134_29 (.A0(\register[2]_c [27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27224), .COUT(n27225), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_29.INIT0 = 16'h5aaa;
    defparam add_134_29.INIT1 = 16'h5aaa;
    defparam add_134_29.INJECT1_0 = "NO";
    defparam add_134_29.INJECT1_1 = "NO";
    CCU2D add_134_27 (.A0(\register[2]_c [25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27223), .COUT(n27224), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_27.INIT0 = 16'h5aaa;
    defparam add_134_27.INIT1 = 16'h5aaa;
    defparam add_134_27.INJECT1_0 = "NO";
    defparam add_134_27.INJECT1_1 = "NO";
    CCU2D add_134_25 (.A0(\register[2]_c [23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27222), .COUT(n27223), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_25.INIT0 = 16'h5aaa;
    defparam add_134_25.INIT1 = 16'h5aaa;
    defparam add_134_25.INJECT1_0 = "NO";
    defparam add_134_25.INJECT1_1 = "NO";
    CCU2D add_134_23 (.A0(\register[2]_c [21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27221), .COUT(n27222), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_23.INIT0 = 16'h5aaa;
    defparam add_134_23.INIT1 = 16'h5aaa;
    defparam add_134_23.INJECT1_0 = "NO";
    defparam add_134_23.INJECT1_1 = "NO";
    FD1P3IX force_pause_151 (.D(\databus[1] ), .SP(n28621), .CD(n33448), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam force_pause_151.GSR = "ENABLED";
    CCU2D add_134_21 (.A0(\register[2]_c [19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27220), .COUT(n27221), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_21.INIT0 = 16'h5aaa;
    defparam add_134_21.INIT1 = 16'h5aaa;
    defparam add_134_21.INJECT1_0 = "NO";
    defparam add_134_21.INJECT1_1 = "NO";
    CCU2D add_134_19 (.A0(\register[2]_c [17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27219), .COUT(n27220), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_19.INIT0 = 16'h5aaa;
    defparam add_134_19.INIT1 = 16'h5aaa;
    defparam add_134_19.INJECT1_0 = "NO";
    defparam add_134_19.INJECT1_1 = "NO";
    CCU2D add_134_17 (.A0(\register[2]_c [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27218), .COUT(n27219), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_17.INIT0 = 16'h5aaa;
    defparam add_134_17.INIT1 = 16'h5aaa;
    defparam add_134_17.INJECT1_0 = "NO";
    defparam add_134_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n31739), .C(\register[2]_c [30]), 
         .D(\register_addr[0] ), .Z(n29504)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0020;
    CCU2D add_134_15 (.A0(\register[2]_c [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27217), .COUT(n27218), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_15.INIT0 = 16'h5aaa;
    defparam add_134_15.INIT1 = 16'h5aaa;
    defparam add_134_15.INJECT1_0 = "NO";
    defparam add_134_15.INJECT1_1 = "NO";
    CCU2D add_134_13 (.A0(\register[2]_c [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27216), .COUT(n27217), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_13.INIT0 = 16'h5aaa;
    defparam add_134_13.INIT1 = 16'h5aaa;
    defparam add_134_13.INJECT1_0 = "NO";
    defparam add_134_13.INJECT1_1 = "NO";
    CCU2D add_134_11 (.A0(\register[2]_c [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27215), .COUT(n27216), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_11.INIT0 = 16'h5aaa;
    defparam add_134_11.INIT1 = 16'h5aaa;
    defparam add_134_11.INJECT1_0 = "NO";
    defparam add_134_11.INJECT1_1 = "NO";
    CCU2D add_134_9 (.A0(\register[2]_c [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27214), .COUT(n27215), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_9.INIT0 = 16'h5aaa;
    defparam add_134_9.INIT1 = 16'h5aaa;
    defparam add_134_9.INJECT1_0 = "NO";
    defparam add_134_9.INJECT1_1 = "NO";
    CCU2D add_134_7 (.A0(\register[2]_c [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27213), .COUT(n27214), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_7.INIT0 = 16'h5aaa;
    defparam add_134_7.INIT1 = 16'h5aaa;
    defparam add_134_7.INJECT1_0 = "NO";
    defparam add_134_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_446 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [31]), .D(\register_addr[0] ), .Z(n29503)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_446.init = 16'h0020;
    CCU2D add_134_5 (.A0(\register[2]_c [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27212), .COUT(n27213), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_5.INIT0 = 16'h5aaa;
    defparam add_134_5.INIT1 = 16'h5aaa;
    defparam add_134_5.INJECT1_0 = "NO";
    defparam add_134_5.INJECT1_1 = "NO";
    CCU2D add_134_3 (.A0(\register[2]_c [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2]_c [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27211), .COUT(n27212), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_3.INIT0 = 16'h5aaa;
    defparam add_134_3.INIT1 = 16'h5aaa;
    defparam add_134_3.INJECT1_0 = "NO";
    defparam add_134_3.INJECT1_1 = "NO";
    CCU2D add_134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27211), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_1.INIT0 = 16'hF000;
    defparam add_134_1.INIT1 = 16'h5555;
    defparam add_134_1.INJECT1_0 = "NO";
    defparam add_134_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_279_4_lut (.A(\register_addr[1] ), .B(n31739), .C(n27707), 
         .D(n31827), .Z(n31702)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_3_lut_rep_279_4_lut.init = 16'h0200;
    LUT4 i2_3_lut_4_lut (.A(\register_addr[1] ), .B(n31739), .C(n14022), 
         .D(\register_addr[0] ), .Z(n9075)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_447 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [29]), .D(\register_addr[0] ), .Z(n29506)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_447.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_448 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [28]), .D(\register_addr[0] ), .Z(n29501)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_448.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_449 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [27]), .D(\register_addr[0] ), .Z(n29505)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_449.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_450 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [26]), .D(\register_addr[0] ), .Z(n29499)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_450.init = 16'h0020;
    LUT4 i1_4_lut (.A(rw), .B(n33447), .C(n29823), .D(\select[1] ), 
         .Z(n28621)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hcdcc;
    LUT4 i1_2_lut_3_lut_4_lut_adj_451 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [25]), .D(\register_addr[0] ), .Z(n29500)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_451.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_452 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [24]), .D(\register_addr[0] ), .Z(n29497)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_452.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_453 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [23]), .D(\register_addr[0] ), .Z(n29486)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_453.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_454 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [22]), .D(\register_addr[0] ), .Z(n29509)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_454.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_455 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [21]), .D(\register_addr[0] ), .Z(n29496)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_455.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_456 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [20]), .D(\register_addr[0] ), .Z(n29491)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_456.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_457 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [19]), .D(\register_addr[0] ), .Z(n29489)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_457.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_458 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [18]), .D(\register_addr[0] ), .Z(n29487)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_458.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_459 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [17]), .D(\register_addr[0] ), .Z(n29507)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_459.init = 16'h0020;
    LUT4 i134_2_lut_rep_408 (.A(prev_clk_1Hz), .B(clk_1Hz), .Z(n31831)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i134_2_lut_rep_408.init = 16'h4444;
    LUT4 i2656_2_lut_3_lut (.A(prev_clk_1Hz), .B(clk_1Hz), .C(n33447), 
         .Z(n9030)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i2656_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_4_lut_adj_460 (.A(\register_addr[0] ), .B(\register[2]_c [3]), 
         .C(n24729), .D(n31720), .Z(n28853)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_460.init = 16'h5450;
    LUT4 i112_2_lut_rep_409 (.A(\register[0] [2]), .B(force_pause), .Z(n31832)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i112_2_lut_rep_409.init = 16'heeee;
    LUT4 i2_3_lut_4_lut_adj_461 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7] ), .D(n27893), .Z(n32)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_461.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_462 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [16]), .D(\register_addr[0] ), .Z(n29495)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_462.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_463 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [15]), .D(\register_addr[0] ), .Z(n29510)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_463.init = 16'h0020;
    LUT4 i2_3_lut_4_lut_adj_464 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_301 ), .D(n27905), .Z(n32_adj_302)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_464.init = 16'h1000;
    LUT4 i15596_2_lut_3_lut_rep_373_4_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(n21959), .D(\register[1][1] ), .Z(n31796)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i15596_2_lut_3_lut_rep_373_4_lut.init = 16'hf0e0;
    LUT4 i14736_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(clk_1Hz), 
         .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i14736_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_465 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [14]), .D(\register_addr[0] ), .Z(n29494)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_465.init = 16'h0020;
    LUT4 i2_3_lut_4_lut_adj_466 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_303 ), .D(n27902), .Z(n32_adj_304)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_466.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_467 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_305 ), .D(n27910), .Z(n34)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_467.init = 16'h1000;
    LUT4 i15592_2_lut_3_lut_rep_374_4_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(n21892), .D(\register[0][1] ), .Z(n31797)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i15592_2_lut_3_lut_rep_374_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_468 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [13]), .D(\register_addr[0] ), .Z(n29508)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_468.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_469 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [12]), .D(\register_addr[0] ), .Z(n29490)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_469.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_470 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [11]), .D(\register_addr[0] ), .Z(n29493)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_470.init = 16'h0020;
    LUT4 i15122_2_lut_rep_375_3_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(\register[0][7] ), .Z(n31798)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i15122_2_lut_rep_375_3_lut.init = 16'h1010;
    LUT4 i23198_2_lut_2_lut_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), 
         .C(n21959), .D(\register[1][1] ), .Z(n21729)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i23198_2_lut_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i23216_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(n31), 
         .D(\state[0] ), .Z(n19)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i23216_3_lut_4_lut.init = 16'h00ef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_471 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [10]), .D(\register_addr[0] ), .Z(n29484)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_471.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_472 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [9]), .D(\register_addr[0] ), .Z(n29483)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_472.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_473 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [8]), .D(\register_addr[0] ), .Z(n29502)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_473.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_474 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [7]), .D(\register_addr[0] ), .Z(n29488)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_474.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_475 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [6]), .D(\register_addr[0] ), .Z(n29485)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_475.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_476 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [5]), .D(\register_addr[0] ), .Z(n29492)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_476.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_477 (.A(\register_addr[1] ), .B(n31739), 
         .C(\register[2]_c [4]), .D(\register_addr[0] ), .Z(n29498)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_477.init = 16'h0020;
    LUT4 i23201_4_lut (.A(\register_addr[2] ), .B(n29738), .C(\register_addr[1] ), 
         .D(\register_addr[0] ), .Z(n29739)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B))) */ ;
    defparam i23201_4_lut.init = 16'h1113;
    LUT4 i28_4_lut (.A(force_pause), .B(\register[2]_c [1]), .C(\register_addr[1] ), 
         .D(\register_addr[0] ), .Z(n21)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i28_4_lut.init = 16'h0fca;
    LUT4 i3_4_lut (.A(n31779), .B(\register_addr[5] ), .C(\register_addr[4] ), 
         .D(n24), .Z(n28729)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut.init = 16'h0100;
    LUT4 i31_4_lut (.A(\register[0] [2]), .B(\register[2]_c [2]), .C(\register_addr[1] ), 
         .D(\register_addr[0] ), .Z(n24)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i31_4_lut.init = 16'h0fca;
    FD1P3AX read_value__i31 (.D(n29503), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29504), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29506), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29501), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29505), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29499), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29500), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29497), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29486), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29509), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29496), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29491), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29489), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29487), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29507), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29495), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29510), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29494), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29508), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29490), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29493), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29484), .SP(n14022), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29483), .SP(n14022), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29502), .SP(n14022), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29488), .SP(n14022), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29485), .SP(n14022), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 i942_3_lut (.A(prev_select), .B(n33447), .C(\select[1] ), .Z(n14022)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(61[5] 104[8])
    defparam i942_3_lut.init = 16'h1010;
    FD1P3AX read_value__i5 (.D(n29492), .SP(n14022), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29498), .SP(n14022), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i4.GSR = "ENABLED";
    LUT4 i114_1_lut (.A(xbee_pause_c), .Z(n178)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(54[26:39])
    defparam i114_1_lut.init = 16'h5555;
    FD1P3IX read_value__i3 (.D(n28853), .SP(n14022), .CD(n9075), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_size_i0_i1 (.D(n29739), .SP(n14022), .CD(n16046), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n31718), .SP(n14022), .CD(n16045), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3AX read_value__i1 (.D(n29452), .SP(n14022), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3AX read_value__i2 (.D(n28729), .SP(n14022), .CK(debug_c_c), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i2.GSR = "ENABLED";
    \ClockDividerP(factor=12000000)  uptime_div (.GND_net(GND_net), .clk_1Hz(clk_1Hz), 
            .debug_c_c(debug_c_c), .n33448(n33448), .n33447(n33447)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(107[28] 109[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (GND_net, clk_1Hz, debug_c_c, 
            n33448, n33447) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output clk_1Hz;
    input debug_c_c;
    input n33448;
    input n33447;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27468;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n27469, n27467, n25, n26, n24, n7589, n27554, n27553, 
        n27552, n27551, n27550, n27549, n27548, n27547, n27546, 
        n27545, n27544, n27543, n2679, n19, n29, n26_adj_562, 
        n32, n30140, n27, n27822, n28, n20, n27482, n27481, 
        n27480, n27479, n27478, n27477, n27476, n27475, n27474, 
        n27473, n27472, n27471, n27470;
    
    CCU2D count_2577_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27468), .COUT(n27469), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_5.INJECT1_0 = "NO";
    defparam count_2577_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27467), .COUT(n27468), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_3.INJECT1_0 = "NO";
    defparam count_2577_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27467), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_1.INIT0 = 16'hF000;
    defparam count_2577_add_4_1.INIT1 = 16'h0555;
    defparam count_2577_add_4_1.INJECT1_0 = "NO";
    defparam count_2577_add_4_1.INJECT1_1 = "NO";
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    FD1S3IX clk_o_14 (.D(n7589), .CK(debug_c_c), .CD(n33448), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D add_20537_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27554), 
          .S0(n7589));
    defparam add_20537_cout.INIT0 = 16'h0000;
    defparam add_20537_cout.INIT1 = 16'h0000;
    defparam add_20537_cout.INJECT1_0 = "NO";
    defparam add_20537_cout.INJECT1_1 = "NO";
    CCU2D add_20537_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27553), .COUT(n27554));
    defparam add_20537_24.INIT0 = 16'h5555;
    defparam add_20537_24.INIT1 = 16'h5555;
    defparam add_20537_24.INJECT1_0 = "NO";
    defparam add_20537_24.INJECT1_1 = "NO";
    CCU2D add_20537_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27552), .COUT(n27553));
    defparam add_20537_22.INIT0 = 16'h5555;
    defparam add_20537_22.INIT1 = 16'h5555;
    defparam add_20537_22.INJECT1_0 = "NO";
    defparam add_20537_22.INJECT1_1 = "NO";
    CCU2D add_20537_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27551), .COUT(n27552));
    defparam add_20537_20.INIT0 = 16'h5555;
    defparam add_20537_20.INIT1 = 16'h5555;
    defparam add_20537_20.INJECT1_0 = "NO";
    defparam add_20537_20.INJECT1_1 = "NO";
    CCU2D add_20537_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27550), .COUT(n27551));
    defparam add_20537_18.INIT0 = 16'h5555;
    defparam add_20537_18.INIT1 = 16'h5555;
    defparam add_20537_18.INJECT1_0 = "NO";
    defparam add_20537_18.INJECT1_1 = "NO";
    CCU2D add_20537_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27549), .COUT(n27550));
    defparam add_20537_16.INIT0 = 16'h5aaa;
    defparam add_20537_16.INIT1 = 16'h5555;
    defparam add_20537_16.INJECT1_0 = "NO";
    defparam add_20537_16.INJECT1_1 = "NO";
    CCU2D add_20537_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27548), .COUT(n27549));
    defparam add_20537_14.INIT0 = 16'h5aaa;
    defparam add_20537_14.INIT1 = 16'h5555;
    defparam add_20537_14.INJECT1_0 = "NO";
    defparam add_20537_14.INJECT1_1 = "NO";
    CCU2D add_20537_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27547), .COUT(n27548));
    defparam add_20537_12.INIT0 = 16'h5555;
    defparam add_20537_12.INIT1 = 16'h5aaa;
    defparam add_20537_12.INJECT1_0 = "NO";
    defparam add_20537_12.INJECT1_1 = "NO";
    CCU2D add_20537_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27546), .COUT(n27547));
    defparam add_20537_10.INIT0 = 16'h5aaa;
    defparam add_20537_10.INIT1 = 16'h5aaa;
    defparam add_20537_10.INJECT1_0 = "NO";
    defparam add_20537_10.INJECT1_1 = "NO";
    CCU2D add_20537_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27545), .COUT(n27546));
    defparam add_20537_8.INIT0 = 16'h5555;
    defparam add_20537_8.INIT1 = 16'h5aaa;
    defparam add_20537_8.INJECT1_0 = "NO";
    defparam add_20537_8.INJECT1_1 = "NO";
    CCU2D add_20537_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27544), .COUT(n27545));
    defparam add_20537_6.INIT0 = 16'h5555;
    defparam add_20537_6.INIT1 = 16'h5555;
    defparam add_20537_6.INJECT1_0 = "NO";
    defparam add_20537_6.INJECT1_1 = "NO";
    CCU2D add_20537_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27543), .COUT(n27544));
    defparam add_20537_4.INIT0 = 16'h5aaa;
    defparam add_20537_4.INIT1 = 16'h5aaa;
    defparam add_20537_4.INJECT1_0 = "NO";
    defparam add_20537_4.INJECT1_1 = "NO";
    CCU2D add_20537_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27543));
    defparam add_20537_2.INIT0 = 16'h7000;
    defparam add_20537_2.INIT1 = 16'h5555;
    defparam add_20537_2.INJECT1_0 = "NO";
    defparam add_20537_2.INJECT1_1 = "NO";
    FD1S3IX count_2577__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2679), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i0.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_562), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i23087_2_lut (.A(n30140), .B(n33447), .Z(n2679)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23087_2_lut.init = 16'heeee;
    LUT4 i23085_4_lut (.A(n27), .B(n27822), .C(n25), .D(n26), .Z(n30140)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i23085_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut_adj_444 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_444.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n27822)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i12_4_lut_adj_445 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_445.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_562)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    FD1S3IX count_2577__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2679), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i1.GSR = "ENABLED";
    FD1S3IX count_2577__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2679), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i2.GSR = "ENABLED";
    FD1S3IX count_2577__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2679), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i3.GSR = "ENABLED";
    FD1S3IX count_2577__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2679), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i4.GSR = "ENABLED";
    FD1S3IX count_2577__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2679), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i5.GSR = "ENABLED";
    FD1S3IX count_2577__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2679), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i6.GSR = "ENABLED";
    FD1S3IX count_2577__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2679), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i7.GSR = "ENABLED";
    FD1S3IX count_2577__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2679), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i8.GSR = "ENABLED";
    FD1S3IX count_2577__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2679), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i9.GSR = "ENABLED";
    FD1S3IX count_2577__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i10.GSR = "ENABLED";
    FD1S3IX count_2577__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i11.GSR = "ENABLED";
    FD1S3IX count_2577__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i12.GSR = "ENABLED";
    FD1S3IX count_2577__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i13.GSR = "ENABLED";
    FD1S3IX count_2577__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i14.GSR = "ENABLED";
    FD1S3IX count_2577__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i15.GSR = "ENABLED";
    FD1S3IX count_2577__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i16.GSR = "ENABLED";
    FD1S3IX count_2577__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i17.GSR = "ENABLED";
    FD1S3IX count_2577__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i18.GSR = "ENABLED";
    FD1S3IX count_2577__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i19.GSR = "ENABLED";
    FD1S3IX count_2577__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i20.GSR = "ENABLED";
    FD1S3IX count_2577__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i21.GSR = "ENABLED";
    FD1S3IX count_2577__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i22.GSR = "ENABLED";
    FD1S3IX count_2577__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i23.GSR = "ENABLED";
    FD1S3IX count_2577__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i24.GSR = "ENABLED";
    FD1S3IX count_2577__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i25.GSR = "ENABLED";
    FD1S3IX count_2577__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i26.GSR = "ENABLED";
    FD1S3IX count_2577__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i27.GSR = "ENABLED";
    FD1S3IX count_2577__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i28.GSR = "ENABLED";
    FD1S3IX count_2577__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i29.GSR = "ENABLED";
    FD1S3IX count_2577__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i30.GSR = "ENABLED";
    FD1S3IX count_2577__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2679), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577__i31.GSR = "ENABLED";
    CCU2D count_2577_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27482), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_33.INIT1 = 16'h0000;
    defparam count_2577_add_4_33.INJECT1_0 = "NO";
    defparam count_2577_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27481), .COUT(n27482), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_31.INJECT1_0 = "NO";
    defparam count_2577_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27480), .COUT(n27481), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_29.INJECT1_0 = "NO";
    defparam count_2577_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27479), .COUT(n27480), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_27.INJECT1_0 = "NO";
    defparam count_2577_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27478), .COUT(n27479), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_25.INJECT1_0 = "NO";
    defparam count_2577_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27477), .COUT(n27478), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_23.INJECT1_0 = "NO";
    defparam count_2577_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27476), .COUT(n27477), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_21.INJECT1_0 = "NO";
    defparam count_2577_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27475), .COUT(n27476), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_19.INJECT1_0 = "NO";
    defparam count_2577_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27474), .COUT(n27475), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_17.INJECT1_0 = "NO";
    defparam count_2577_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27473), .COUT(n27474), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_15.INJECT1_0 = "NO";
    defparam count_2577_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27472), .COUT(n27473), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_13.INJECT1_0 = "NO";
    defparam count_2577_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27471), .COUT(n27472), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_11.INJECT1_0 = "NO";
    defparam count_2577_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27470), .COUT(n27471), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_9.INJECT1_0 = "NO";
    defparam count_2577_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2577_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27469), .COUT(n27470), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2577_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2577_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2577_add_4_7.INJECT1_0 = "NO";
    defparam count_2577_add_4_7.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (read_value, debug_c_c, n2669, 
            n9093, n33450, VCC_net, GND_net, Stepper_A_nFault_c, \read_size[0] , 
            n8940, Stepper_A_M0_c_0, n14252, n579, prev_select, n31741, 
            n33447, \register_addr[1] , Stepper_A_M1_c_1, n32, n32_adj_294, 
            prev_step_clk, step_clk, n31711, n22, n32_adj_295, prev_step_clk_adj_296, 
            step_clk_adj_297, n31712, \register_addr[0] , n22_adj_298, 
            prev_step_clk_adj_299, n34, step_clk_adj_300, n31713, n24, 
            n33446, n191, n185, n33448, n33449, n33451, \read_size[2] , 
            n29590, n31700, n33453, databus, Stepper_A_M2_c_2, Stepper_A_Dir_c, 
            Stepper_A_En_c, \control_reg[7] , n8885, n31784, n27905, 
            n3700, limit_c_3, Stepper_A_Step_c, n8261) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2669;
    input n9093;
    input n33450;
    input VCC_net;
    input GND_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n8940;
    output Stepper_A_M0_c_0;
    input n14252;
    input n579;
    output prev_select;
    input n31741;
    input n33447;
    input \register_addr[1] ;
    output Stepper_A_M1_c_1;
    input n32;
    input n32_adj_294;
    input prev_step_clk;
    input step_clk;
    output n31711;
    output n22;
    input n32_adj_295;
    input prev_step_clk_adj_296;
    input step_clk_adj_297;
    output n31712;
    input \register_addr[0] ;
    output n22_adj_298;
    input prev_step_clk_adj_299;
    input n34;
    input step_clk_adj_300;
    output n31713;
    output n24;
    input n33446;
    input n191;
    output n185;
    input n33448;
    input n33449;
    input n33451;
    output \read_size[2] ;
    input n29590;
    input n31700;
    input n33453;
    input [31:0]databus;
    output Stepper_A_M2_c_2;
    output Stepper_A_Dir_c;
    output Stepper_A_En_c;
    output \control_reg[7] ;
    input n8885;
    input n31784;
    output n27905;
    input n3700;
    input limit_c_3;
    output Stepper_A_Step_c;
    input n8261;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30088;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n3701;
    
    wire fault_latched, prev_step_clk_c, step_clk_c, limit_latched, 
        n182, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n14292;
    wire [31:0]n100;
    
    wire n11687, n16, n30046, n31896, n31895, n31894, n31710, 
        n22_c, n27330;
    wire [31:0]n224;
    
    wire n27329, n27328, n27327, n27326, n27325, n27324, n27323, 
        n30086, n27322, n27321, n27320, n27319, n30087, n27318, 
        n27317, n27316, n27315, int_step, n30044, n30045;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n49, n62_adj_553, n58_adj_554, n50_adj_555, n41, n60_adj_556, 
        n54_adj_557, n42_adj_558, n52_adj_559, n38_adj_560, n56, n46_adj_561;
    wire [7:0]n8260;
    wire [31:0]n7150;
    
    FD1P3IX read_value__i0 (.D(n30088), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3701[0]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n8940), .SP(n2669), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n14252), .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk_c), .CK(debug_c_c), .Q(prev_step_clk_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n14292), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31741), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i5286_3_lut (.A(prev_limit_latched), .B(n33447), .C(limit_latched), 
         .Z(n11687)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i5286_3_lut.init = 16'hdcdc;
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n16), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30046), .SP(n2669), .CD(n9093), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3AX read_value__i1 (.D(n31896), .SP(n2669), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 n30089_bdd_4_lut_then_4_lut (.A(steps_reg[1]), .B(fault_latched), 
         .C(n9093), .D(\register_addr[1] ), .Z(n31895)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam n30089_bdd_4_lut_then_4_lut.init = 16'h0a0c;
    LUT4 n30089_bdd_4_lut_else_4_lut (.A(Stepper_A_M1_c_1), .B(n9093), .C(div_factor_reg[1]), 
         .D(\register_addr[1] ), .Z(n31894)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam n30089_bdd_4_lut_else_4_lut.init = 16'h3022;
    LUT4 i2_3_lut_rep_287 (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .Z(n31710)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_287.init = 16'h2020;
    LUT4 i1_4_lut_4_lut (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .D(n33447), .Z(n22_c)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut.init = 16'h002c;
    LUT4 i2_3_lut_rep_288 (.A(n32_adj_294), .B(prev_step_clk), .C(step_clk), 
         .Z(n31711)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_288.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_adj_440 (.A(n32_adj_294), .B(prev_step_clk), .C(step_clk), 
         .D(n33447), .Z(n22)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_440.init = 16'h002c;
    LUT4 i2_3_lut_rep_289 (.A(n32_adj_295), .B(prev_step_clk_adj_296), .C(step_clk_adj_297), 
         .Z(n31712)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_289.init = 16'h2020;
    LUT4 i14808_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14808_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_4_lut_adj_441 (.A(n32_adj_295), .B(prev_step_clk_adj_296), 
         .C(step_clk_adj_297), .D(n33447), .Z(n22_adj_298)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_441.init = 16'h002c;
    LUT4 i2_3_lut_rep_290 (.A(prev_step_clk_adj_299), .B(n34), .C(step_clk_adj_300), 
         .Z(n31713)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_290.init = 16'h4040;
    LUT4 i14809_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14809_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_4_lut_adj_442 (.A(prev_step_clk_adj_299), .B(n34), .C(step_clk_adj_300), 
         .D(n33447), .Z(n24)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_442.init = 16'h004a;
    LUT4 i14810_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14810_4_lut.init = 16'hc088;
    LUT4 i14811_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14811_4_lut.init = 16'hc088;
    LUT4 i14812_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14812_4_lut.init = 16'hc088;
    LUT4 i14813_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14813_4_lut.init = 16'hc088;
    LUT4 i14814_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14814_4_lut.init = 16'hc088;
    LUT4 i14815_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14815_4_lut.init = 16'hc088;
    LUT4 i14816_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14816_4_lut.init = 16'hc088;
    LUT4 i14817_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14817_4_lut.init = 16'hc088;
    LUT4 i14818_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14818_4_lut.init = 16'hc088;
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[20]), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n16)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i14819_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14819_4_lut.init = 16'hc088;
    LUT4 i14820_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14820_4_lut.init = 16'hc088;
    LUT4 i14821_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14821_4_lut.init = 16'hc088;
    LUT4 i2_3_lut_4_lut (.A(n31741), .B(prev_select), .C(n33446), .D(n191), 
         .Z(n185)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_4_lut.init = 16'h0200;
    LUT4 i14822_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14822_4_lut.init = 16'hc088;
    LUT4 i14823_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14823_4_lut.init = 16'hc088;
    LUT4 i14824_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14824_4_lut.init = 16'hc088;
    LUT4 i14825_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14825_4_lut.init = 16'hc088;
    LUT4 i14826_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14826_4_lut.init = 16'hc088;
    LUT4 i14827_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14827_4_lut.init = 16'hc088;
    LUT4 i14828_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14828_4_lut.init = 16'hc088;
    LUT4 i14829_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14829_4_lut.init = 16'hc088;
    LUT4 i14830_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14830_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27330), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27329), .COUT(n27330), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27328), .COUT(n27329), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27327), .COUT(n27328), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27326), .COUT(n27327), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27325), .COUT(n27326), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27324), .COUT(n27325), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27323), .COUT(n27324), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    LUT4 i22933_3_lut (.A(Stepper_A_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22933_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27322), .COUT(n27323), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27321), .COUT(n27322), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27320), .COUT(n27321), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27319), .COUT(n27320), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    LUT4 i22934_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22934_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27318), .COUT(n27319), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27317), .COUT(n27318), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27316), .COUT(n27317), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27315), .COUT(n27316), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk_c), .D1(prev_step_clk_c), 
          .COUT(n27315), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    FD1P3AX int_step_182 (.D(n31710), .SP(n22_c), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3701[31]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3701[30]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3701[29]), .CK(debug_c_c), .CD(n33449), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3701[28]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3701[27]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3701[26]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3701[25]), .CK(debug_c_c), .CD(n33449), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3701[24]), .CK(debug_c_c), .CD(n33449), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3701[23]), .CK(debug_c_c), .CD(n33449), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3701[22]), .CK(debug_c_c), .CD(n33449), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3701[21]), .CK(debug_c_c), .CD(n33449), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3701[20]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3701[19]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3701[18]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3701[17]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3701[16]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3701[15]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3701[14]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3701[13]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3701[12]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3701[11]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3701[10]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3701[9]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3701[8]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3701[7]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3701[6]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3701[5]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3701[4]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3701[3]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3701[2]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3701[1]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    PFUMX i22893 (.BLUT(n30044), .ALUT(n30045), .C0(\register_addr[0] ), 
          .Z(n30046));
    FD1P3AX read_size__i2 (.D(n29590), .SP(n2669), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n31700), .PD(n33453), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n31700), .CD(n33453), 
            .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n31700), .PD(n33453), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n31700), .CD(n33453), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n31700), .PD(n33453), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n31700), .PD(n33453), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n31700), .CD(n11687), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n8885), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n8885), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n8885), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n8885), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n8885), .PD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n8885), .PD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n8885), .PD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n8885), .PD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n8885), .PD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n8885), .PD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n8885), .PD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n8885), .CD(n31784), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=603, LSE_RLINE=616 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_553), .C(n58_adj_554), .D(n50_adj_555), 
         .Z(n27905)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[20]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_556), .C(n54_adj_557), .D(n42_adj_558), 
         .Z(n62_adj_553)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52_adj_559), .C(n38_adj_560), 
         .D(steps_reg[24]), .Z(n58_adj_554)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50_adj_555)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[25]), .B(steps_reg[26]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[9]), .B(n56), .C(n46_adj_561), .D(steps_reg[2]), 
         .Z(n60_adj_556)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[16]), .B(steps_reg[22]), .C(steps_reg[4]), 
         .D(steps_reg[18]), .Z(n54_adj_557)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[29]), .B(steps_reg[0]), .Z(n42_adj_558)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[17]), .B(steps_reg[3]), .C(steps_reg[6]), 
         .D(steps_reg[10]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[12]), .Z(n46_adj_561)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[28]), .B(steps_reg[7]), .C(steps_reg[30]), 
         .D(steps_reg[8]), .Z(n52_adj_559)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[1]), .B(steps_reg[13]), .Z(n38_adj_560)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    PFUMX i22935 (.BLUT(n30086), .ALUT(n30087), .C0(\register_addr[1] ), 
          .Z(n30088));
    LUT4 i14834_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8260[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14834_2_lut.init = 16'h2222;
    LUT4 mux_1947_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7150[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1947_i4_3_lut.init = 16'hcaca;
    LUT4 i14833_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8260[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14833_2_lut.init = 16'h2222;
    LUT4 mux_1947_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7150[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1947_i5_3_lut.init = 16'hcaca;
    LUT4 i14832_2_lut (.A(Stepper_A_Dir_c), .B(\register_addr[0] ), .Z(n8260[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14832_2_lut.init = 16'h2222;
    LUT4 mux_1947_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7150[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1947_i6_3_lut.init = 16'hcaca;
    LUT4 i14831_2_lut (.A(Stepper_A_En_c), .B(\register_addr[0] ), .Z(n8260[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14831_2_lut.init = 16'h2222;
    LUT4 mux_1947_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7150[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1947_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1947_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n7150[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1947_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3700), 
         .Z(n3701[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3700), 
         .Z(n3701[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3700), 
         .Z(n3701[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3700), 
         .Z(n3701[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3700), 
         .Z(n3701[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3700), 
         .Z(n3701[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3700), 
         .Z(n3701[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3700), 
         .Z(n3701[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3700), 
         .Z(n3701[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3700), 
         .Z(n3701[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3700), 
         .Z(n3701[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3700), 
         .Z(n3701[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3700), 
         .Z(n3701[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3700), 
         .Z(n3701[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i19_3_lut.init = 16'hcaca;
    LUT4 i22891_3_lut (.A(Stepper_A_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22891_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3700), 
         .Z(n3701[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3700), 
         .Z(n3701[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3700), 
         .Z(n3701[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3700), 
         .Z(n3701[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3700), 
         .Z(n3701[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3700), 
         .Z(n3701[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3700), 
         .Z(n3701[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3700), 
         .Z(n3701[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3700), .Z(n3701[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i10_3_lut.init = 16'hcaca;
    LUT4 i22892_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22892_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3700), .Z(n3701[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3700), .Z(n3701[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3700), .Z(n3701[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3700), .Z(n3701[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3700), .Z(n3701[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3700), .Z(n3701[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3700), .Z(n3701[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3700), .Z(n3701[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1499_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3700), .Z(n3701[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1499_i1_3_lut.init = 16'hcaca;
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(n8885), .B(n33447), .Z(n14292)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_443 (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_443.init = 16'h9999;
    PFUMX mux_1951_i4 (.BLUT(n8260[3]), .ALUT(n7150[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_1951_i5 (.BLUT(n8260[4]), .ALUT(n7150[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX i23760 (.BLUT(n31894), .ALUT(n31895), .C0(\register_addr[0] ), 
          .Z(n31896));
    PFUMX mux_1951_i6 (.BLUT(n8260[5]), .ALUT(n7150[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1951_i7 (.BLUT(n8260[6]), .ALUT(n7150[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    PFUMX mux_1951_i8 (.BLUT(n8261), .ALUT(n7150[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    ClockDivider_U9 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk_c), 
            .debug_c_c(debug_c_c), .n33448(n33448), .n33447(n33447), .div_factor_reg({div_factor_reg})) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (GND_net, step_clk, debug_c_c, n33448, n33447, 
            div_factor_reg) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n33448;
    input n33447;
    input [31:0]div_factor_reg;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27257;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n27258, n27466;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27256, n27465, n27464, n27255, n27463, n27254, n27462, 
        n27461, n27460, n27459, n27458, n27253, n27457, n27456, 
        n27455, n27454, n27453, n27252, n27452, n27451, n27251, 
        n7936, n27066, n7971, n31691, n27065, n27064, n27063, 
        n27062, n27061, n27060, n27059, n27058, n27057, n27056, 
        n27055, n27054, n27053, n27052, n27051, n27050, n27049, 
        n27048, n27047, n27046, n27045, n27044, n27043, n27042, 
        n27041, n27040, n27039, n27038, n27037, n27036, n27035, 
        n27034, n8005, n27033, n27032, n27031, n27030, n27029, 
        n27028, n27027, n27026, n27025, n27024, n27023, n27022, 
        n27021, n27020, n27019, n16112, n27266, n27265, n27264, 
        n27263, n27262, n27261, n27260, n27259;
    
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27257), .COUT(n27258), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27466), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_33.INIT1 = 16'h0000;
    defparam count_2581_add_4_33.INJECT1_0 = "NO";
    defparam count_2581_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27256), .COUT(n27257), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27465), .COUT(n27466), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_31.INJECT1_0 = "NO";
    defparam count_2581_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27464), .COUT(n27465), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_29.INJECT1_0 = "NO";
    defparam count_2581_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27255), .COUT(n27256), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27463), .COUT(n27464), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_27.INJECT1_0 = "NO";
    defparam count_2581_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27254), .COUT(n27255), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27462), .COUT(n27463), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_25.INJECT1_0 = "NO";
    defparam count_2581_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27461), .COUT(n27462), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_23.INJECT1_0 = "NO";
    defparam count_2581_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27460), .COUT(n27461), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_21.INJECT1_0 = "NO";
    defparam count_2581_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27459), .COUT(n27460), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_19.INJECT1_0 = "NO";
    defparam count_2581_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27458), .COUT(n27459), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_17.INJECT1_0 = "NO";
    defparam count_2581_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27253), .COUT(n27254), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27457), .COUT(n27458), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_15.INJECT1_0 = "NO";
    defparam count_2581_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27456), .COUT(n27457), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_13.INJECT1_0 = "NO";
    defparam count_2581_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27455), .COUT(n27456), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_11.INJECT1_0 = "NO";
    defparam count_2581_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27454), .COUT(n27455), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_9.INJECT1_0 = "NO";
    defparam count_2581_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27453), .COUT(n27454), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_7.INJECT1_0 = "NO";
    defparam count_2581_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27252), .COUT(n27253), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27452), .COUT(n27453), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_5.INJECT1_0 = "NO";
    defparam count_2581_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27451), .COUT(n27452), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2581_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2581_add_4_3.INJECT1_0 = "NO";
    defparam count_2581_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2581_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27451), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581_add_4_1.INIT0 = 16'hF000;
    defparam count_2581_add_4_1.INIT1 = 16'h0555;
    defparam count_2581_add_4_1.INJECT1_0 = "NO";
    defparam count_2581_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27251), .COUT(n27252), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27251), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7936), .CK(debug_c_c), .CD(n33448), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2009_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27066), .S1(n7936));
    defparam sub_2009_add_2_33.INIT0 = 16'h5555;
    defparam sub_2009_add_2_33.INIT1 = 16'h0000;
    defparam sub_2009_add_2_33.INJECT1_0 = "NO";
    defparam sub_2009_add_2_33.INJECT1_1 = "NO";
    LUT4 i1013_2_lut_rep_268 (.A(n7971), .B(n33447), .Z(n31691)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1013_2_lut_rep_268.init = 16'heeee;
    CCU2D sub_2009_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27065), .COUT(n27066));
    defparam sub_2009_add_2_31.INIT0 = 16'h5999;
    defparam sub_2009_add_2_31.INIT1 = 16'h5999;
    defparam sub_2009_add_2_31.INJECT1_0 = "NO";
    defparam sub_2009_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27064), .COUT(n27065));
    defparam sub_2009_add_2_29.INIT0 = 16'h5999;
    defparam sub_2009_add_2_29.INIT1 = 16'h5999;
    defparam sub_2009_add_2_29.INJECT1_0 = "NO";
    defparam sub_2009_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27063), .COUT(n27064));
    defparam sub_2009_add_2_27.INIT0 = 16'h5999;
    defparam sub_2009_add_2_27.INIT1 = 16'h5999;
    defparam sub_2009_add_2_27.INJECT1_0 = "NO";
    defparam sub_2009_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27062), .COUT(n27063));
    defparam sub_2009_add_2_25.INIT0 = 16'h5999;
    defparam sub_2009_add_2_25.INIT1 = 16'h5999;
    defparam sub_2009_add_2_25.INJECT1_0 = "NO";
    defparam sub_2009_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27061), .COUT(n27062));
    defparam sub_2009_add_2_23.INIT0 = 16'h5999;
    defparam sub_2009_add_2_23.INIT1 = 16'h5999;
    defparam sub_2009_add_2_23.INJECT1_0 = "NO";
    defparam sub_2009_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27060), .COUT(n27061));
    defparam sub_2009_add_2_21.INIT0 = 16'h5999;
    defparam sub_2009_add_2_21.INIT1 = 16'h5999;
    defparam sub_2009_add_2_21.INJECT1_0 = "NO";
    defparam sub_2009_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27059), .COUT(n27060));
    defparam sub_2009_add_2_19.INIT0 = 16'h5999;
    defparam sub_2009_add_2_19.INIT1 = 16'h5999;
    defparam sub_2009_add_2_19.INJECT1_0 = "NO";
    defparam sub_2009_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27058), .COUT(n27059));
    defparam sub_2009_add_2_17.INIT0 = 16'h5999;
    defparam sub_2009_add_2_17.INIT1 = 16'h5999;
    defparam sub_2009_add_2_17.INJECT1_0 = "NO";
    defparam sub_2009_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27057), .COUT(n27058));
    defparam sub_2009_add_2_15.INIT0 = 16'h5999;
    defparam sub_2009_add_2_15.INIT1 = 16'h5999;
    defparam sub_2009_add_2_15.INJECT1_0 = "NO";
    defparam sub_2009_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27056), .COUT(n27057));
    defparam sub_2009_add_2_13.INIT0 = 16'h5999;
    defparam sub_2009_add_2_13.INIT1 = 16'h5999;
    defparam sub_2009_add_2_13.INJECT1_0 = "NO";
    defparam sub_2009_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27055), .COUT(n27056));
    defparam sub_2009_add_2_11.INIT0 = 16'h5999;
    defparam sub_2009_add_2_11.INIT1 = 16'h5999;
    defparam sub_2009_add_2_11.INJECT1_0 = "NO";
    defparam sub_2009_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27054), .COUT(n27055));
    defparam sub_2009_add_2_9.INIT0 = 16'h5999;
    defparam sub_2009_add_2_9.INIT1 = 16'h5999;
    defparam sub_2009_add_2_9.INJECT1_0 = "NO";
    defparam sub_2009_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27053), .COUT(n27054));
    defparam sub_2009_add_2_7.INIT0 = 16'h5999;
    defparam sub_2009_add_2_7.INIT1 = 16'h5999;
    defparam sub_2009_add_2_7.INJECT1_0 = "NO";
    defparam sub_2009_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27052), .COUT(n27053));
    defparam sub_2009_add_2_5.INIT0 = 16'h5999;
    defparam sub_2009_add_2_5.INIT1 = 16'h5999;
    defparam sub_2009_add_2_5.INJECT1_0 = "NO";
    defparam sub_2009_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27051), .COUT(n27052));
    defparam sub_2009_add_2_3.INIT0 = 16'h5999;
    defparam sub_2009_add_2_3.INIT1 = 16'h5999;
    defparam sub_2009_add_2_3.INJECT1_0 = "NO";
    defparam sub_2009_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2009_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27051));
    defparam sub_2009_add_2_1.INIT0 = 16'h0000;
    defparam sub_2009_add_2_1.INIT1 = 16'h5999;
    defparam sub_2009_add_2_1.INJECT1_0 = "NO";
    defparam sub_2009_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27050), .S1(n7971));
    defparam sub_2011_add_2_33.INIT0 = 16'h5999;
    defparam sub_2011_add_2_33.INIT1 = 16'h0000;
    defparam sub_2011_add_2_33.INJECT1_0 = "NO";
    defparam sub_2011_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27049), .COUT(n27050));
    defparam sub_2011_add_2_31.INIT0 = 16'h5999;
    defparam sub_2011_add_2_31.INIT1 = 16'h5999;
    defparam sub_2011_add_2_31.INJECT1_0 = "NO";
    defparam sub_2011_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27048), .COUT(n27049));
    defparam sub_2011_add_2_29.INIT0 = 16'h5999;
    defparam sub_2011_add_2_29.INIT1 = 16'h5999;
    defparam sub_2011_add_2_29.INJECT1_0 = "NO";
    defparam sub_2011_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27047), .COUT(n27048));
    defparam sub_2011_add_2_27.INIT0 = 16'h5999;
    defparam sub_2011_add_2_27.INIT1 = 16'h5999;
    defparam sub_2011_add_2_27.INJECT1_0 = "NO";
    defparam sub_2011_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27046), .COUT(n27047));
    defparam sub_2011_add_2_25.INIT0 = 16'h5999;
    defparam sub_2011_add_2_25.INIT1 = 16'h5999;
    defparam sub_2011_add_2_25.INJECT1_0 = "NO";
    defparam sub_2011_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27045), .COUT(n27046));
    defparam sub_2011_add_2_23.INIT0 = 16'h5999;
    defparam sub_2011_add_2_23.INIT1 = 16'h5999;
    defparam sub_2011_add_2_23.INJECT1_0 = "NO";
    defparam sub_2011_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27044), .COUT(n27045));
    defparam sub_2011_add_2_21.INIT0 = 16'h5999;
    defparam sub_2011_add_2_21.INIT1 = 16'h5999;
    defparam sub_2011_add_2_21.INJECT1_0 = "NO";
    defparam sub_2011_add_2_21.INJECT1_1 = "NO";
    FD1S3IX count_2581__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i0.GSR = "ENABLED";
    CCU2D sub_2011_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27043), .COUT(n27044));
    defparam sub_2011_add_2_19.INIT0 = 16'h5999;
    defparam sub_2011_add_2_19.INIT1 = 16'h5999;
    defparam sub_2011_add_2_19.INJECT1_0 = "NO";
    defparam sub_2011_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27042), .COUT(n27043));
    defparam sub_2011_add_2_17.INIT0 = 16'h5999;
    defparam sub_2011_add_2_17.INIT1 = 16'h5999;
    defparam sub_2011_add_2_17.INJECT1_0 = "NO";
    defparam sub_2011_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27041), .COUT(n27042));
    defparam sub_2011_add_2_15.INIT0 = 16'h5999;
    defparam sub_2011_add_2_15.INIT1 = 16'h5999;
    defparam sub_2011_add_2_15.INJECT1_0 = "NO";
    defparam sub_2011_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27040), .COUT(n27041));
    defparam sub_2011_add_2_13.INIT0 = 16'h5999;
    defparam sub_2011_add_2_13.INIT1 = 16'h5999;
    defparam sub_2011_add_2_13.INJECT1_0 = "NO";
    defparam sub_2011_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27039), .COUT(n27040));
    defparam sub_2011_add_2_11.INIT0 = 16'h5999;
    defparam sub_2011_add_2_11.INIT1 = 16'h5999;
    defparam sub_2011_add_2_11.INJECT1_0 = "NO";
    defparam sub_2011_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27038), .COUT(n27039));
    defparam sub_2011_add_2_9.INIT0 = 16'h5999;
    defparam sub_2011_add_2_9.INIT1 = 16'h5999;
    defparam sub_2011_add_2_9.INJECT1_0 = "NO";
    defparam sub_2011_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27037), .COUT(n27038));
    defparam sub_2011_add_2_7.INIT0 = 16'h5999;
    defparam sub_2011_add_2_7.INIT1 = 16'h5999;
    defparam sub_2011_add_2_7.INJECT1_0 = "NO";
    defparam sub_2011_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27036), .COUT(n27037));
    defparam sub_2011_add_2_5.INIT0 = 16'h5999;
    defparam sub_2011_add_2_5.INIT1 = 16'h5999;
    defparam sub_2011_add_2_5.INJECT1_0 = "NO";
    defparam sub_2011_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27035), .COUT(n27036));
    defparam sub_2011_add_2_3.INIT0 = 16'h5999;
    defparam sub_2011_add_2_3.INIT1 = 16'h5999;
    defparam sub_2011_add_2_3.INJECT1_0 = "NO";
    defparam sub_2011_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2011_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27035));
    defparam sub_2011_add_2_1.INIT0 = 16'h0000;
    defparam sub_2011_add_2_1.INIT1 = 16'h5999;
    defparam sub_2011_add_2_1.INJECT1_0 = "NO";
    defparam sub_2011_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27034), .S1(n8005));
    defparam sub_2012_add_2_33.INIT0 = 16'hf555;
    defparam sub_2012_add_2_33.INIT1 = 16'h0000;
    defparam sub_2012_add_2_33.INJECT1_0 = "NO";
    defparam sub_2012_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27033), .COUT(n27034));
    defparam sub_2012_add_2_31.INIT0 = 16'hf555;
    defparam sub_2012_add_2_31.INIT1 = 16'hf555;
    defparam sub_2012_add_2_31.INJECT1_0 = "NO";
    defparam sub_2012_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27032), .COUT(n27033));
    defparam sub_2012_add_2_29.INIT0 = 16'hf555;
    defparam sub_2012_add_2_29.INIT1 = 16'hf555;
    defparam sub_2012_add_2_29.INJECT1_0 = "NO";
    defparam sub_2012_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27031), .COUT(n27032));
    defparam sub_2012_add_2_27.INIT0 = 16'hf555;
    defparam sub_2012_add_2_27.INIT1 = 16'hf555;
    defparam sub_2012_add_2_27.INJECT1_0 = "NO";
    defparam sub_2012_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27030), .COUT(n27031));
    defparam sub_2012_add_2_25.INIT0 = 16'hf555;
    defparam sub_2012_add_2_25.INIT1 = 16'hf555;
    defparam sub_2012_add_2_25.INJECT1_0 = "NO";
    defparam sub_2012_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27029), .COUT(n27030));
    defparam sub_2012_add_2_23.INIT0 = 16'hf555;
    defparam sub_2012_add_2_23.INIT1 = 16'hf555;
    defparam sub_2012_add_2_23.INJECT1_0 = "NO";
    defparam sub_2012_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27028), .COUT(n27029));
    defparam sub_2012_add_2_21.INIT0 = 16'hf555;
    defparam sub_2012_add_2_21.INIT1 = 16'hf555;
    defparam sub_2012_add_2_21.INJECT1_0 = "NO";
    defparam sub_2012_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27027), .COUT(n27028));
    defparam sub_2012_add_2_19.INIT0 = 16'hf555;
    defparam sub_2012_add_2_19.INIT1 = 16'hf555;
    defparam sub_2012_add_2_19.INJECT1_0 = "NO";
    defparam sub_2012_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27026), .COUT(n27027));
    defparam sub_2012_add_2_17.INIT0 = 16'hf555;
    defparam sub_2012_add_2_17.INIT1 = 16'hf555;
    defparam sub_2012_add_2_17.INJECT1_0 = "NO";
    defparam sub_2012_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27025), .COUT(n27026));
    defparam sub_2012_add_2_15.INIT0 = 16'hf555;
    defparam sub_2012_add_2_15.INIT1 = 16'hf555;
    defparam sub_2012_add_2_15.INJECT1_0 = "NO";
    defparam sub_2012_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27024), .COUT(n27025));
    defparam sub_2012_add_2_13.INIT0 = 16'hf555;
    defparam sub_2012_add_2_13.INIT1 = 16'hf555;
    defparam sub_2012_add_2_13.INJECT1_0 = "NO";
    defparam sub_2012_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27023), .COUT(n27024));
    defparam sub_2012_add_2_11.INIT0 = 16'hf555;
    defparam sub_2012_add_2_11.INIT1 = 16'hf555;
    defparam sub_2012_add_2_11.INJECT1_0 = "NO";
    defparam sub_2012_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27022), .COUT(n27023));
    defparam sub_2012_add_2_9.INIT0 = 16'hf555;
    defparam sub_2012_add_2_9.INIT1 = 16'hf555;
    defparam sub_2012_add_2_9.INJECT1_0 = "NO";
    defparam sub_2012_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27021), .COUT(n27022));
    defparam sub_2012_add_2_7.INIT0 = 16'hf555;
    defparam sub_2012_add_2_7.INIT1 = 16'hf555;
    defparam sub_2012_add_2_7.INJECT1_0 = "NO";
    defparam sub_2012_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27020), .COUT(n27021));
    defparam sub_2012_add_2_5.INIT0 = 16'hf555;
    defparam sub_2012_add_2_5.INIT1 = 16'hf555;
    defparam sub_2012_add_2_5.INJECT1_0 = "NO";
    defparam sub_2012_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2012_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27019), .COUT(n27020));
    defparam sub_2012_add_2_3.INIT0 = 16'hf555;
    defparam sub_2012_add_2_3.INIT1 = 16'hf555;
    defparam sub_2012_add_2_3.INJECT1_0 = "NO";
    defparam sub_2012_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    CCU2D sub_2012_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27019));
    defparam sub_2012_add_2_1.INIT0 = 16'h0000;
    defparam sub_2012_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2012_add_2_1.INJECT1_0 = "NO";
    defparam sub_2012_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31691), .PD(n16112), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1S3IX count_2581__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i1.GSR = "ENABLED";
    FD1S3IX count_2581__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i2.GSR = "ENABLED";
    FD1S3IX count_2581__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i3.GSR = "ENABLED";
    FD1S3IX count_2581__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i4.GSR = "ENABLED";
    FD1S3IX count_2581__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i5.GSR = "ENABLED";
    FD1S3IX count_2581__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i6.GSR = "ENABLED";
    FD1S3IX count_2581__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i7.GSR = "ENABLED";
    FD1S3IX count_2581__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i8.GSR = "ENABLED";
    FD1S3IX count_2581__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i9.GSR = "ENABLED";
    FD1S3IX count_2581__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i10.GSR = "ENABLED";
    FD1S3IX count_2581__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i11.GSR = "ENABLED";
    FD1S3IX count_2581__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i12.GSR = "ENABLED";
    FD1S3IX count_2581__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i13.GSR = "ENABLED";
    FD1S3IX count_2581__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i14.GSR = "ENABLED";
    FD1S3IX count_2581__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i15.GSR = "ENABLED";
    FD1S3IX count_2581__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i16.GSR = "ENABLED";
    FD1S3IX count_2581__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i17.GSR = "ENABLED";
    FD1S3IX count_2581__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i18.GSR = "ENABLED";
    FD1S3IX count_2581__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i19.GSR = "ENABLED";
    FD1S3IX count_2581__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i20.GSR = "ENABLED";
    FD1S3IX count_2581__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i21.GSR = "ENABLED";
    FD1S3IX count_2581__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i22.GSR = "ENABLED";
    FD1S3IX count_2581__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i23.GSR = "ENABLED";
    FD1S3IX count_2581__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i24.GSR = "ENABLED";
    FD1S3IX count_2581__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i25.GSR = "ENABLED";
    FD1S3IX count_2581__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i26.GSR = "ENABLED";
    FD1S3IX count_2581__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i27.GSR = "ENABLED";
    FD1S3IX count_2581__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i28.GSR = "ENABLED";
    FD1S3IX count_2581__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i29.GSR = "ENABLED";
    FD1S3IX count_2581__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i30.GSR = "ENABLED";
    FD1S3IX count_2581__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31691), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2581__i31.GSR = "ENABLED";
    LUT4 i9706_2_lut_3_lut (.A(n7971), .B(n33447), .C(n8005), .Z(n16112)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9706_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27266), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27265), .COUT(n27266), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27264), .COUT(n27265), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27263), .COUT(n27264), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27262), .COUT(n27263), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27261), .COUT(n27262), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27260), .COUT(n27261), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27259), .COUT(n27260), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27258), .COUT(n27259), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31691), .CD(n16112), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP_SP(factor=12000000) 
//

module \ClockDividerP_SP(factor=12000000)  (GND_net, clk_10Hz, debug_c_c, 
            n33448, n33447) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output clk_10Hz;
    input debug_c_c;
    input n33448;
    input n33447;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(86[13:18])
    
    wire n27, n29, n26, n32, n28, n26_adj_540, n20, n28_adj_541, 
        n24, n16, n27450;
    wire [31:0]n134;
    
    wire n27449, n27448, n27447, n27446, n27445, n27444, n27443, 
        n31790, n27442, n27441, n27440, n27439, n27438, n27437, 
        n27436, n27435, n28242, n2672, n30143, n29996, n30029, 
        n29994, n29992, n29998;
    
    LUT4 i10_4_lut (.A(count[12]), .B(count[20]), .C(count[18]), .D(count[23]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(n29), .B(count[4]), .C(n26), .D(count[16]), .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[11]), .B(count[6]), .C(count[21]), .D(count[9]), 
         .Z(n28)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i12_4_lut (.A(count[17]), .B(count[7]), .C(count[0]), .D(count[5]), 
         .Z(n29)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i9_3_lut (.A(count[2]), .B(count[1]), .C(count[3]), .Z(n26)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i9_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(count[19]), .B(n26_adj_540), .C(n20), .D(count[26]), 
         .Z(n28_adj_541)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[10]), .B(count[30]), .C(count[8]), .D(count[14]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[31]), .B(count[22]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i11_4_lut_adj_439 (.A(count[27]), .B(count[13]), .C(count[29]), 
         .D(count[25]), .Z(n26_adj_540)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i11_4_lut_adj_439.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[28]), .B(count[24]), .Z(n20)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i5_2_lut.init = 16'heeee;
    CCU2D count_2576_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27450), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_33.INIT1 = 16'h0000;
    defparam count_2576_add_4_33.INJECT1_0 = "NO";
    defparam count_2576_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27449), .COUT(n27450), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_31.INJECT1_0 = "NO";
    defparam count_2576_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27448), .COUT(n27449), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_29.INJECT1_0 = "NO";
    defparam count_2576_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27447), .COUT(n27448), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_27.INJECT1_0 = "NO";
    defparam count_2576_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27446), .COUT(n27447), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_25.INJECT1_0 = "NO";
    defparam count_2576_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27445), .COUT(n27446), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_23.INJECT1_0 = "NO";
    defparam count_2576_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27444), .COUT(n27445), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_21.INJECT1_0 = "NO";
    defparam count_2576_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27443), .COUT(n27444), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_19.INJECT1_0 = "NO";
    defparam count_2576_add_4_19.INJECT1_1 = "NO";
    LUT4 i14_4_lut_rep_367 (.A(count[15]), .B(n28_adj_541), .C(n24), .D(n16), 
         .Z(n31790)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i14_4_lut_rep_367.init = 16'hfffe;
    CCU2D count_2576_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27442), .COUT(n27443), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_17.INJECT1_0 = "NO";
    defparam count_2576_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27441), .COUT(n27442), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_15.INJECT1_0 = "NO";
    defparam count_2576_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27440), .COUT(n27441), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_13.INJECT1_0 = "NO";
    defparam count_2576_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27439), .COUT(n27440), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_11.INJECT1_0 = "NO";
    defparam count_2576_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27438), .COUT(n27439), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_9.INJECT1_0 = "NO";
    defparam count_2576_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27437), .COUT(n27438), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_7.INJECT1_0 = "NO";
    defparam count_2576_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27436), .COUT(n27437), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_5.INJECT1_0 = "NO";
    defparam count_2576_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27435), .COUT(n27436), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2576_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2576_add_4_3.INJECT1_0 = "NO";
    defparam count_2576_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2576_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27435), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576_add_4_1.INIT0 = 16'hF000;
    defparam count_2576_add_4_1.INIT1 = 16'h0555;
    defparam count_2576_add_4_1.INJECT1_0 = "NO";
    defparam count_2576_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_13 (.D(n28242), .CK(debug_c_c), .CD(n33448), .Q(clk_10Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(88[9] 107[6])
    defparam clk_o_13.GSR = "ENABLED";
    FD1S3IX count_2576__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2672), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i0.GSR = "ENABLED";
    LUT4 i23090_2_lut (.A(n30143), .B(n33447), .Z(n2672)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23090_2_lut.init = 16'heeee;
    LUT4 i23088_4_lut (.A(n31790), .B(n29996), .C(n30029), .D(n29994), 
         .Z(n30143)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i23088_4_lut.init = 16'h4000;
    LUT4 i22844_4_lut (.A(count[18]), .B(count[2]), .C(count[1]), .D(count[11]), 
         .Z(n29996)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22844_4_lut.init = 16'h8000;
    LUT4 i22876_4_lut (.A(n29992), .B(count[9]), .C(n29998), .D(count[0]), 
         .Z(n30029)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22876_4_lut.init = 16'h8000;
    LUT4 i22842_4_lut (.A(count[3]), .B(count[12]), .C(count[5]), .D(count[17]), 
         .Z(n29994)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22842_4_lut.init = 16'h8000;
    LUT4 i22840_4_lut (.A(count[20]), .B(count[7]), .C(count[23]), .D(count[21]), 
         .Z(n29992)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22840_4_lut.init = 16'h8000;
    LUT4 i22846_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n29998)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22846_3_lut.init = 16'h8080;
    FD1S3IX count_2576__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2672), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i1.GSR = "ENABLED";
    FD1S3IX count_2576__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2672), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i2.GSR = "ENABLED";
    FD1S3IX count_2576__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2672), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i3.GSR = "ENABLED";
    FD1S3IX count_2576__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2672), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i4.GSR = "ENABLED";
    FD1S3IX count_2576__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2672), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i5.GSR = "ENABLED";
    FD1S3IX count_2576__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2672), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i6.GSR = "ENABLED";
    FD1S3IX count_2576__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2672), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i7.GSR = "ENABLED";
    FD1S3IX count_2576__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2672), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i8.GSR = "ENABLED";
    FD1S3IX count_2576__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2672), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i9.GSR = "ENABLED";
    FD1S3IX count_2576__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i10.GSR = "ENABLED";
    FD1S3IX count_2576__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i11.GSR = "ENABLED";
    FD1S3IX count_2576__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i12.GSR = "ENABLED";
    FD1S3IX count_2576__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i13.GSR = "ENABLED";
    FD1S3IX count_2576__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i14.GSR = "ENABLED";
    FD1S3IX count_2576__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i15.GSR = "ENABLED";
    FD1S3IX count_2576__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i16.GSR = "ENABLED";
    FD1S3IX count_2576__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i17.GSR = "ENABLED";
    FD1S3IX count_2576__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i18.GSR = "ENABLED";
    FD1S3IX count_2576__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i19.GSR = "ENABLED";
    FD1S3IX count_2576__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i20.GSR = "ENABLED";
    FD1S3IX count_2576__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i21.GSR = "ENABLED";
    FD1S3IX count_2576__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i22.GSR = "ENABLED";
    FD1S3IX count_2576__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i23.GSR = "ENABLED";
    FD1S3IX count_2576__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i24.GSR = "ENABLED";
    FD1S3IX count_2576__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i25.GSR = "ENABLED";
    FD1S3IX count_2576__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i26.GSR = "ENABLED";
    FD1S3IX count_2576__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i27.GSR = "ENABLED";
    FD1S3IX count_2576__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i28.GSR = "ENABLED";
    FD1S3IX count_2576__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i29.GSR = "ENABLED";
    FD1S3IX count_2576__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i30.GSR = "ENABLED";
    FD1S3IX count_2576__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2672), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2576__i31.GSR = "ENABLED";
    LUT4 i23154_4_lut_4_lut (.A(n31790), .B(n28), .C(n32), .D(n27), 
         .Z(n28242)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i23154_4_lut_4_lut.init = 16'h0001;
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (\read_value[18] , read_value, n31719, n47, \read_value[18]_adj_91 , 
            n6, n31703, databus_out, rw, \read_value[18]_adj_92 , 
            read_value_adj_293, n31716, n46, n3, databus, \read_value[17]_adj_125 , 
            \read_value[17]_adj_126 , n6_adj_127, \read_value[6]_adj_128 , 
            n31733, n33446, \read_value[17]_adj_129 , \read_value[6]_adj_130 , 
            n3_adj_131, \select[7] , \read_value[16]_adj_132 , \read_value[16]_adj_133 , 
            n6_adj_134, \read_value[16]_adj_135 , n3_adj_136, \read_value[15]_adj_137 , 
            \read_value[15]_adj_138 , n6_adj_139, \read_value[15]_adj_140 , 
            \register_addr[0] , n8, \read_value[7]_adj_141 , n3_adj_142, 
            \read_value[14]_adj_143 , \read_value[14]_adj_144 , n6_adj_145, 
            n8_adj_146, \read_value[14]_adj_147 , n3_adj_148, \read_value[13]_adj_149 , 
            \read_value[13]_adj_150 , n6_adj_151, \read_value[13]_adj_152 , 
            \read_value[7]_adj_153 , n3_adj_154, n3_adj_155, \read_value[31]_adj_156 , 
            \read_value[12]_adj_157 , \read_value[12]_adj_158 , n6_adj_159, 
            \read_value[31]_adj_160 , n6_adj_161, \read_value[12]_adj_162 , 
            \read_value[31]_adj_163 , n3_adj_164, \read_value[11]_adj_165 , 
            \read_value[11]_adj_166 , n6_adj_167, \read_value[11]_adj_168 , 
            \register_addr[2] , \register_addr[1] , n3_adj_169, \read_value[10]_adj_170 , 
            \read_value[10]_adj_171 , n6_adj_172, n3_adj_173, \read_value[30]_adj_174 , 
            \read_value[30]_adj_175 , n6_adj_176, \read_value[10]_adj_177 , 
            \read_value[30]_adj_178 , n3_adj_179, \read_value[29]_adj_180 , 
            \read_value[29]_adj_181 , n6_adj_182, \read_value[29]_adj_183 , 
            n3_adj_184, \read_value[9]_adj_185 , n3_adj_186, \read_value[28]_adj_187 , 
            \read_value[9]_adj_188 , n6_adj_189, \read_value[28]_adj_190 , 
            n6_adj_191, \read_value[28]_adj_192 , \read_value[9]_adj_193 , 
            n3_adj_194, \read_value[27]_adj_195 , n3_adj_196, \read_value[27]_adj_197 , 
            n6_adj_198, \read_value[27]_adj_199 , \read_value[8]_adj_200 , 
            \read_value[8]_adj_201 , n6_adj_202, \read_value[8]_adj_203 , 
            n3_adj_204, \read_value[26]_adj_205 , \read_value[26]_adj_206 , 
            n6_adj_207, \read_value[26]_adj_208 , n3_adj_209, \read_value[25]_adj_210 , 
            \read_value[25]_adj_211 , n6_adj_212, \read_value[25]_adj_213 , 
            \read_size[0] , \read_size[0]_adj_214 , \select[2] , n31780, 
            n9, n29694, n14, n3_adj_215, \select[4] , \read_size[0]_adj_216 , 
            n55, n31762, n10, read_size, n31732, \select[1] , \read_size[0]_adj_218 , 
            n31741, n6_adj_219, \read_size[2]_adj_220 , \reg_size[2] , 
            n9_adj_221, \read_size[2]_adj_222 , \read_value[24]_adj_223 , 
            \read_value[24]_adj_224 , n6_adj_225, \read_size[2]_adj_226 , 
            n2, \read_value[5]_adj_227 , n5, n8_adj_228, \read_value[24]_adj_229 , 
            n3_adj_230, \read_value[23]_adj_231 , \read_value[23]_adj_232 , 
            n6_adj_233, n2_adj_234, \read_value[23]_adj_235 , \read_value[5]_adj_236 , 
            \read_value[6]_adj_237 , n5_adj_238, n3_adj_239, \read_value[5]_adj_240 , 
            \read_value[22]_adj_241 , \read_value[22]_adj_242 , n6_adj_243, 
            \read_value[22]_adj_244 , n3_adj_245, \read_value[21]_adj_246 , 
            \read_value[21]_adj_247 , n6_adj_248, \read_value[21]_adj_249 , 
            n3_adj_250, n31841, \sendcount[1] , n12795, \read_value[20]_adj_251 , 
            \read_value[20]_adj_252 , n6_adj_253, \read_value[20]_adj_254 , 
            n2_adj_255, n3_adj_256, \read_value[19]_adj_257 , \read_value[19]_adj_258 , 
            n6_adj_259, \read_value[4]_adj_260 , n5_adj_261, n8_adj_262, 
            \read_value[19]_adj_263 , n3_adj_264, n8_adj_265, \read_value[4]_adj_266 , 
            \read_value[4]_adj_267 , n2_adj_268, \read_value[3]_adj_269 , 
            n5_adj_270, n8_adj_271, \read_value[3]_adj_272 , \read_value[3]_adj_273 , 
            \read_value[7]_adj_274 , n5_adj_275, n29738, n2_adj_276, 
            \read_value[2]_adj_277 , n5_adj_278, n8_adj_279, \read_value[2]_adj_280 , 
            \read_value[2]_adj_281 , n1, n5_adj_282, \read_value[0]_adj_283 , 
            n2_adj_284, \read_value[0]_adj_285 , \read_value[1]_adj_286 , 
            n4, n2_adj_287, \read_value[1]_adj_288 , n31746, n2_adj_289, 
            \read_value[0]_adj_290 , n5_adj_291, GND_net, debug_c_c, 
            n31694, rc_ch8_c, n27918, n30160, n30216, n13719, rc_ch7_c, 
            n27933, n30195, n14176, n30205, rc_ch4_c, n27937, n30182, 
            n14182, n30191, n30197, rc_ch3_c, n27924, n14183, n30189, 
            n30186, rc_ch2_c, n27915, n14186, n30218, n29930, n14187, 
            n9_adj_292, rc_ch1_c, n30152, n30184, n27912) /* synthesis syn_module_defined=1 */ ;
    input \read_value[18] ;
    input [31:0]read_value;
    input n31719;
    input n47;
    input \read_value[18]_adj_91 ;
    input n6;
    input n31703;
    input [31:0]databus_out;
    input rw;
    input \read_value[18]_adj_92 ;
    input [31:0]read_value_adj_293;
    input n31716;
    input n46;
    input n3;
    output [31:0]databus;
    input \read_value[17]_adj_125 ;
    input \read_value[17]_adj_126 ;
    input n6_adj_127;
    input \read_value[6]_adj_128 ;
    input n31733;
    input n33446;
    input \read_value[17]_adj_129 ;
    input \read_value[6]_adj_130 ;
    input n3_adj_131;
    input \select[7] ;
    input \read_value[16]_adj_132 ;
    input \read_value[16]_adj_133 ;
    input n6_adj_134;
    input \read_value[16]_adj_135 ;
    input n3_adj_136;
    input \read_value[15]_adj_137 ;
    input \read_value[15]_adj_138 ;
    input n6_adj_139;
    input \read_value[15]_adj_140 ;
    input \register_addr[0] ;
    input n8;
    input \read_value[7]_adj_141 ;
    input n3_adj_142;
    input \read_value[14]_adj_143 ;
    input \read_value[14]_adj_144 ;
    input n6_adj_145;
    input n8_adj_146;
    input \read_value[14]_adj_147 ;
    input n3_adj_148;
    input \read_value[13]_adj_149 ;
    input \read_value[13]_adj_150 ;
    input n6_adj_151;
    input \read_value[13]_adj_152 ;
    input \read_value[7]_adj_153 ;
    input n3_adj_154;
    input n3_adj_155;
    input \read_value[31]_adj_156 ;
    input \read_value[12]_adj_157 ;
    input \read_value[12]_adj_158 ;
    input n6_adj_159;
    input \read_value[31]_adj_160 ;
    input n6_adj_161;
    input \read_value[12]_adj_162 ;
    input \read_value[31]_adj_163 ;
    input n3_adj_164;
    input \read_value[11]_adj_165 ;
    input \read_value[11]_adj_166 ;
    input n6_adj_167;
    input \read_value[11]_adj_168 ;
    input \register_addr[2] ;
    input \register_addr[1] ;
    input n3_adj_169;
    input \read_value[10]_adj_170 ;
    input \read_value[10]_adj_171 ;
    input n6_adj_172;
    input n3_adj_173;
    input \read_value[30]_adj_174 ;
    input \read_value[30]_adj_175 ;
    input n6_adj_176;
    input \read_value[10]_adj_177 ;
    input \read_value[30]_adj_178 ;
    input n3_adj_179;
    input \read_value[29]_adj_180 ;
    input \read_value[29]_adj_181 ;
    input n6_adj_182;
    input \read_value[29]_adj_183 ;
    input n3_adj_184;
    input \read_value[9]_adj_185 ;
    input n3_adj_186;
    input \read_value[28]_adj_187 ;
    input \read_value[9]_adj_188 ;
    input n6_adj_189;
    input \read_value[28]_adj_190 ;
    input n6_adj_191;
    input \read_value[28]_adj_192 ;
    input \read_value[9]_adj_193 ;
    input n3_adj_194;
    input \read_value[27]_adj_195 ;
    input n3_adj_196;
    input \read_value[27]_adj_197 ;
    input n6_adj_198;
    input \read_value[27]_adj_199 ;
    input \read_value[8]_adj_200 ;
    input \read_value[8]_adj_201 ;
    input n6_adj_202;
    input \read_value[8]_adj_203 ;
    input n3_adj_204;
    input \read_value[26]_adj_205 ;
    input \read_value[26]_adj_206 ;
    input n6_adj_207;
    input \read_value[26]_adj_208 ;
    input n3_adj_209;
    input \read_value[25]_adj_210 ;
    input \read_value[25]_adj_211 ;
    input n6_adj_212;
    input \read_value[25]_adj_213 ;
    input \read_size[0] ;
    input \read_size[0]_adj_214 ;
    input \select[2] ;
    input n31780;
    output n9;
    input n29694;
    output n14;
    input n3_adj_215;
    input \select[4] ;
    input \read_size[0]_adj_216 ;
    input n55;
    input n31762;
    output n10;
    input [2:0]read_size;
    input n31732;
    input \select[1] ;
    input \read_size[0]_adj_218 ;
    input n31741;
    input n6_adj_219;
    input \read_size[2]_adj_220 ;
    output \reg_size[2] ;
    input n9_adj_221;
    input \read_size[2]_adj_222 ;
    input \read_value[24]_adj_223 ;
    input \read_value[24]_adj_224 ;
    input n6_adj_225;
    input \read_size[2]_adj_226 ;
    input n2;
    input \read_value[5]_adj_227 ;
    input n5;
    input n8_adj_228;
    input \read_value[24]_adj_229 ;
    input n3_adj_230;
    input \read_value[23]_adj_231 ;
    input \read_value[23]_adj_232 ;
    input n6_adj_233;
    input n2_adj_234;
    input \read_value[23]_adj_235 ;
    input \read_value[5]_adj_236 ;
    input \read_value[6]_adj_237 ;
    input n5_adj_238;
    input n3_adj_239;
    input \read_value[5]_adj_240 ;
    input \read_value[22]_adj_241 ;
    input \read_value[22]_adj_242 ;
    input n6_adj_243;
    input \read_value[22]_adj_244 ;
    input n3_adj_245;
    input \read_value[21]_adj_246 ;
    input \read_value[21]_adj_247 ;
    input n6_adj_248;
    input \read_value[21]_adj_249 ;
    input n3_adj_250;
    output n31841;
    input \sendcount[1] ;
    output n12795;
    input \read_value[20]_adj_251 ;
    input \read_value[20]_adj_252 ;
    input n6_adj_253;
    input \read_value[20]_adj_254 ;
    input n2_adj_255;
    input n3_adj_256;
    input \read_value[19]_adj_257 ;
    input \read_value[19]_adj_258 ;
    input n6_adj_259;
    input \read_value[4]_adj_260 ;
    input n5_adj_261;
    input n8_adj_262;
    input \read_value[19]_adj_263 ;
    input n3_adj_264;
    input n8_adj_265;
    input \read_value[4]_adj_266 ;
    input \read_value[4]_adj_267 ;
    input n2_adj_268;
    input \read_value[3]_adj_269 ;
    input n5_adj_270;
    input n8_adj_271;
    input \read_value[3]_adj_272 ;
    input \read_value[3]_adj_273 ;
    input \read_value[7]_adj_274 ;
    input n5_adj_275;
    input n29738;
    input n2_adj_276;
    input \read_value[2]_adj_277 ;
    input n5_adj_278;
    input n8_adj_279;
    input \read_value[2]_adj_280 ;
    input \read_value[2]_adj_281 ;
    input n1;
    input n5_adj_282;
    input \read_value[0]_adj_283 ;
    input n2_adj_284;
    input \read_value[0]_adj_285 ;
    input \read_value[1]_adj_286 ;
    input n4;
    input n2_adj_287;
    input \read_value[1]_adj_288 ;
    input n31746;
    input n2_adj_289;
    input \read_value[0]_adj_290 ;
    input n5_adj_291;
    input GND_net;
    input debug_c_c;
    input n31694;
    input rc_ch8_c;
    input n27918;
    output n30160;
    output n30216;
    input n13719;
    input rc_ch7_c;
    input n27933;
    output n30195;
    input n14176;
    output n30205;
    input rc_ch4_c;
    input n27937;
    output n30182;
    input n14182;
    output n30191;
    output n30197;
    input rc_ch3_c;
    input n27924;
    input n14183;
    output n30189;
    output n30186;
    input rc_ch2_c;
    input n27915;
    input n14186;
    output n30218;
    output n29930;
    input n14187;
    input n9_adj_292;
    input rc_ch1_c;
    output n30152;
    output n30184;
    input n27912;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire n31780 /* synthesis SET_AS_NETWORK=n31780 */ ;
    wire n31762 /* synthesis SET_AS_NETWORK=n31762 */ ;
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n9_c, n12, n14_c, n5_c, n9_adj_195, n14_adj_196, n5_adj_197, 
        n12_adj_200, n14_adj_203;
    wire [7:0]read_value_adj_538;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(210[12:22])
    
    wire n46_adj_208, n12_adj_209, n9_adj_210, n14_adj_211, n5_adj_213;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(211[12:21])
    
    wire n176, n12_adj_216, n9_adj_220, n14_adj_221, n5_adj_223, n12_adj_226;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31558, n12_adj_230, n16, n14_adj_233, n9_adj_234, n14_adj_235, 
        n5_adj_237, n12_adj_240, n12_adj_242, n16_adj_244;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31098, n9_adj_247, n14_adj_248, n5_adj_250, n31096, n12_adj_253;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31095, n1030;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31099, n9_adj_259, n14_adj_260, n5_adj_262, n9_adj_263, 
        n14_adj_264, n5_adj_266, n12_adj_270, n30707, n12_adj_273, 
        n30708, n31557, n31560, n30710, n985, n31561, n9_adj_279, 
        n14_adj_280, n5_adj_282_c, n30711, n12_adj_285, n30842, n30839, 
        n30843, n30841, n30840, n9_adj_289, n14_adj_290, n5_adj_292, 
        n12_adj_295, n9_adj_297, n14_adj_298, n5_adj_300, n31205, 
        n12_adj_303, n31206, n31208, n1000, n31209, n9_adj_309, 
        n14_adj_310, n5_adj_312, n31228, n31229, n12_adj_315, n9_adj_319, 
        n14_adj_320, n5_adj_322, n31231, n9_adj_324, n14_adj_325, 
        n5_adj_327, n12_adj_330, n1045, n31232, n12_adj_333, n9_adj_339, 
        n14_adj_340, n5_adj_342, n9_adj_344, n14_adj_345, n5_adj_347, 
        n12_adj_349, n12_adj_355, n9_adj_359, n14_adj_360, n5_adj_362, 
        n31243, n31242, n12_adj_365, n30838, n30837, n9_adj_369, 
        n14_adj_370, n5_adj_372, n12_adj_375, n31245, n31246, n30712, 
        n30709, n30713, n31271, n1060, n31272, n12_adj_382, n9_adj_384, 
        n14_adj_385, n5_adj_387, n10_adj_391, n8_adj_393, n31269, 
        n12_adj_398, n17, n6_adj_402, n16_adj_403, n31268, n14_adj_404, 
        n31744, n31211, n31101, n31248, n31234, n31274, n12_adj_408, 
        n9_adj_412, n14_adj_413, n5_adj_415, n12_adj_418, n17_adj_420, 
        n6_adj_421, n16_adj_422, n9_adj_430, n14_adj_431, n5_adj_433, 
        n12_adj_437, n1015, n9_adj_441, n14_adj_442, n5_adj_444, n12_adj_447, 
        n9_adj_451, n14_adj_452, n5_adj_454, n12_adj_457, n31562, 
        n31559, n31563, n17_adj_461, n6_adj_462, n16_adj_463, n9_adj_465, 
        n14_adj_466, n5_adj_468, n12_adj_471, n14_adj_474, n12_adj_482, 
        n17_adj_487, n6_adj_488, n16_adj_489, n14_adj_492, n12_adj_495, 
        n6_adj_501, n17_adj_504, n31273, n31270, n17_adj_505, n6_adj_506, 
        n16_adj_507, n31247, n31244, n14_adj_510, n12_adj_513, n31233, 
        n31230, n18, n14_adj_518, n31210, n31207, n16_adj_522, n14_adj_526, 
        n11, n31100, n31097, n17_adj_531, n6_adj_532;
    
    LUT4 i1_4_lut (.A(\read_value[18] ), .B(read_value[18]), .C(n31719), 
         .D(n47), .Z(n9_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i6_4_lut (.A(\read_value[18]_adj_91 ), .B(n12), .C(n6), .D(n31703), 
         .Z(n14_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 Select_4160_i5_2_lut (.A(databus_out[18]), .B(rw), .Z(n5_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4160_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut (.A(\read_value[18]_adj_92 ), .B(read_value_adj_293[18]), 
         .C(n31716), .D(n46), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut.init = 16'heca0;
    LUT4 i7_4_lut (.A(n9_adj_195), .B(n14_adj_196), .C(n3), .D(n5_adj_197), 
         .Z(databus[17])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_304 (.A(\read_value[17]_adj_125 ), .B(read_value[17]), 
         .C(n31719), .D(n47), .Z(n9_adj_195)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_304.init = 16'heca0;
    LUT4 i6_4_lut_adj_305 (.A(\read_value[17]_adj_126 ), .B(n12_adj_200), 
         .C(n6_adj_127), .D(n31703), .Z(n14_adj_196)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_305.init = 16'hfefc;
    LUT4 i4_4_lut_adj_306 (.A(read_value_adj_293[6]), .B(\read_value[6]_adj_128 ), 
         .C(n46), .D(n31733), .Z(n14_adj_203)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_306.init = 16'heca0;
    LUT4 Select_4163_i5_2_lut (.A(databus_out[17]), .B(n33446), .Z(n5_adj_197)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4163_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_307 (.A(\read_value[17]_adj_129 ), .B(read_value_adj_293[17]), 
         .C(n31716), .D(n46), .Z(n12_adj_200)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_307.init = 16'heca0;
    LUT4 i2_4_lut (.A(\read_value[6]_adj_130 ), .B(read_value_adj_538[6]), 
         .C(n31703), .D(n46_adj_208), .Z(n12_adj_209)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 i7_4_lut_adj_308 (.A(n9_adj_210), .B(n14_adj_211), .C(n3_adj_131), 
         .D(n5_adj_213), .Z(databus[16])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_308.init = 16'hfffe;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_309 (.A(\read_value[16]_adj_132 ), .B(read_value[16]), 
         .C(n31719), .D(n47), .Z(n9_adj_210)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_309.init = 16'heca0;
    LUT4 i6_4_lut_adj_310 (.A(\read_value[16]_adj_133 ), .B(n12_adj_216), 
         .C(n6_adj_134), .D(n31703), .Z(n14_adj_211)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_310.init = 16'hfefc;
    LUT4 Select_4166_i5_2_lut (.A(databus_out[16]), .B(rw), .Z(n5_adj_213)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4166_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_311 (.A(\read_value[16]_adj_135 ), .B(read_value_adj_293[16]), 
         .C(n31716), .D(n46), .Z(n12_adj_216)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_311.init = 16'heca0;
    LUT4 i7_4_lut_adj_312 (.A(n9_adj_220), .B(n14_adj_221), .C(n3_adj_136), 
         .D(n5_adj_223), .Z(databus[15])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_312.init = 16'hfffe;
    LUT4 i1_4_lut_adj_313 (.A(\read_value[15]_adj_137 ), .B(read_value[15]), 
         .C(n31719), .D(n47), .Z(n9_adj_220)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_313.init = 16'heca0;
    LUT4 i6_4_lut_adj_314 (.A(\read_value[15]_adj_138 ), .B(n12_adj_226), 
         .C(n6_adj_139), .D(n31703), .Z(n14_adj_221)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_314.init = 16'hfefc;
    LUT4 Select_4169_i5_2_lut (.A(databus_out[15]), .B(rw), .Z(n5_adj_223)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4169_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_315 (.A(\read_value[15]_adj_140 ), .B(read_value_adj_293[15]), 
         .C(n31716), .D(n46), .Z(n12_adj_226)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_315.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23725 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n31558)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23725.init = 16'he4e4;
    LUT4 i6_4_lut_adj_316 (.A(read_value[7]), .B(n12_adj_230), .C(n8), 
         .D(n47), .Z(n16)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_316.init = 16'hfefc;
    LUT4 i4_4_lut_adj_317 (.A(read_value_adj_293[7]), .B(\read_value[7]_adj_141 ), 
         .C(n46), .D(n31733), .Z(n14_adj_233)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_317.init = 16'heca0;
    LUT4 i7_4_lut_adj_318 (.A(n9_adj_234), .B(n14_adj_235), .C(n3_adj_142), 
         .D(n5_adj_237), .Z(databus[14])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_318.init = 16'hfffe;
    LUT4 i1_4_lut_adj_319 (.A(\read_value[14]_adj_143 ), .B(read_value[14]), 
         .C(n31719), .D(n47), .Z(n9_adj_234)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_319.init = 16'heca0;
    LUT4 i6_4_lut_adj_320 (.A(\read_value[14]_adj_144 ), .B(n12_adj_240), 
         .C(n6_adj_145), .D(n31703), .Z(n14_adj_235)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_320.init = 16'hfefc;
    LUT4 i6_4_lut_adj_321 (.A(read_value[0]), .B(n12_adj_242), .C(n8_adj_146), 
         .D(n47), .Z(n16_adj_244)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_321.init = 16'hfefc;
    LUT4 Select_4172_i5_2_lut (.A(databus_out[14]), .B(rw), .Z(n5_adj_237)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4172_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_322 (.A(\read_value[14]_adj_147 ), .B(read_value_adj_293[14]), 
         .C(n31716), .D(n46), .Z(n12_adj_240)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_322.init = 16'heca0;
    LUT4 n1030_bdd_3_lut_23496 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n31098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1030_bdd_3_lut_23496.init = 16'hcaca;
    LUT4 i7_4_lut_adj_323 (.A(n9_adj_247), .B(n14_adj_248), .C(n3_adj_148), 
         .D(n5_adj_250), .Z(databus[13])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_323.init = 16'hfffe;
    LUT4 i1_4_lut_adj_324 (.A(\read_value[13]_adj_149 ), .B(read_value[13]), 
         .C(n31719), .D(n47), .Z(n9_adj_247)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_324.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23512 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n31096)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23512.init = 16'he4e4;
    LUT4 i6_4_lut_adj_325 (.A(\read_value[13]_adj_150 ), .B(n12_adj_253), 
         .C(n6_adj_151), .D(n31703), .Z(n14_adj_248)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_325.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_23511 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n31095)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23511.init = 16'h2222;
    LUT4 n1030_bdd_3_lut_23733 (.A(n1030), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n31099)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1030_bdd_3_lut_23733.init = 16'he2e2;
    LUT4 Select_4175_i5_2_lut (.A(databus_out[13]), .B(rw), .Z(n5_adj_250)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4175_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_326 (.A(\read_value[13]_adj_152 ), .B(read_value_adj_293[13]), 
         .C(n31716), .D(n46), .Z(n12_adj_253)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_326.init = 16'heca0;
    LUT4 i2_4_lut_adj_327 (.A(\read_value[7]_adj_153 ), .B(read_value_adj_538[7]), 
         .C(n31703), .D(n46_adj_208), .Z(n12_adj_230)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_327.init = 16'heca0;
    LUT4 i7_4_lut_adj_328 (.A(n9_adj_259), .B(n14_adj_260), .C(n3_adj_154), 
         .D(n5_adj_262), .Z(databus[12])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_328.init = 16'hfffe;
    LUT4 i7_4_lut_adj_329 (.A(n9_adj_263), .B(n14_adj_264), .C(n3_adj_155), 
         .D(n5_adj_266), .Z(databus[31])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_329.init = 16'hfffe;
    LUT4 i1_4_lut_adj_330 (.A(\read_value[31]_adj_156 ), .B(read_value[31]), 
         .C(n31719), .D(n47), .Z(n9_adj_263)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_330.init = 16'heca0;
    LUT4 i1_4_lut_adj_331 (.A(\read_value[12]_adj_157 ), .B(read_value[12]), 
         .C(n31719), .D(n47), .Z(n9_adj_259)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_331.init = 16'heca0;
    LUT4 i6_4_lut_adj_332 (.A(\read_value[12]_adj_158 ), .B(n12_adj_270), 
         .C(n6_adj_159), .D(n31703), .Z(n14_adj_260)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_332.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_23407 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n30707)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23407.init = 16'h2222;
    LUT4 i6_4_lut_adj_333 (.A(\read_value[31]_adj_160 ), .B(n12_adj_273), 
         .C(n6_adj_161), .D(n31703), .Z(n14_adj_264)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_333.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_23408 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n30708)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23408.init = 16'he4e4;
    LUT4 Select_4121_i5_2_lut (.A(databus_out[31]), .B(rw), .Z(n5_adj_266)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4121_i5_2_lut.init = 16'h2222;
    LUT4 Select_4178_i5_2_lut (.A(databus_out[12]), .B(rw), .Z(n5_adj_262)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4178_i5_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_2_lut_23724 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n31557)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23724.init = 16'h2222;
    LUT4 i4_4_lut_adj_334 (.A(\read_value[12]_adj_162 ), .B(read_value_adj_293[12]), 
         .C(n31716), .D(n46), .Z(n12_adj_270)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_334.init = 16'heca0;
    LUT4 n985_bdd_3_lut_23681 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n31560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n985_bdd_3_lut_23681.init = 16'hcaca;
    LUT4 \register_1[[4__bdd_3_lut_23471  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n30710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_23471 .init = 16'hcaca;
    LUT4 i4_4_lut_adj_335 (.A(\read_value[31]_adj_163 ), .B(read_value_adj_293[31]), 
         .C(n31716), .D(n46), .Z(n12_adj_273)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_335.init = 16'heca0;
    LUT4 n985_bdd_3_lut_23927 (.A(n985), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n31561)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n985_bdd_3_lut_23927.init = 16'he2e2;
    LUT4 i7_4_lut_adj_336 (.A(n9_adj_279), .B(n14_adj_280), .C(n3_adj_164), 
         .D(n5_adj_282_c), .Z(databus[11])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_336.init = 16'hfffe;
    LUT4 i1_4_lut_adj_337 (.A(\read_value[11]_adj_165 ), .B(read_value[11]), 
         .C(n31719), .D(n47), .Z(n9_adj_279)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_337.init = 16'heca0;
    LUT4 \register_1[[4__bdd_2_lut_23472  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n30711)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_23472 .init = 16'h8888;
    LUT4 i6_4_lut_adj_338 (.A(\read_value[11]_adj_166 ), .B(n12_adj_285), 
         .C(n6_adj_167), .D(n31703), .Z(n14_adj_280)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_338.init = 16'hfefc;
    LUT4 Select_4181_i5_2_lut (.A(databus_out[11]), .B(rw), .Z(n5_adj_282_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4181_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_339 (.A(\read_value[11]_adj_168 ), .B(read_value_adj_293[11]), 
         .C(n31716), .D(n46), .Z(n12_adj_285)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_339.init = 16'heca0;
    L6MUX21 i23414 (.D0(n30842), .D1(n30839), .SD(\register_addr[2] ), 
            .Z(n30843));
    PFUMX i23412 (.BLUT(n30841), .ALUT(n30840), .C0(\register_addr[1] ), 
          .Z(n30842));
    LUT4 i7_4_lut_adj_340 (.A(n9_adj_289), .B(n14_adj_290), .C(n3_adj_169), 
         .D(n5_adj_292), .Z(databus[10])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_340.init = 16'hfffe;
    LUT4 i1_4_lut_adj_341 (.A(\read_value[10]_adj_170 ), .B(read_value[10]), 
         .C(n31719), .D(n47), .Z(n9_adj_289)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_341.init = 16'heca0;
    LUT4 i6_4_lut_adj_342 (.A(\read_value[10]_adj_171 ), .B(n12_adj_295), 
         .C(n6_adj_172), .D(n31703), .Z(n14_adj_290)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_342.init = 16'hfefc;
    LUT4 i7_4_lut_adj_343 (.A(n9_adj_297), .B(n14_adj_298), .C(n3_adj_173), 
         .D(n5_adj_300), .Z(databus[30])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_343.init = 16'hfffe;
    LUT4 register_addr_1__bdd_2_lut_23552 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n31205)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23552.init = 16'h2222;
    LUT4 i1_4_lut_adj_344 (.A(\read_value[30]_adj_174 ), .B(read_value[30]), 
         .C(n31719), .D(n47), .Z(n9_adj_297)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_344.init = 16'heca0;
    LUT4 i6_4_lut_adj_345 (.A(\read_value[30]_adj_175 ), .B(n12_adj_303), 
         .C(n6_adj_176), .D(n31703), .Z(n14_adj_298)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_345.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_23553 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n31206)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23553.init = 16'he4e4;
    LUT4 n1000_bdd_3_lut_23538 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n31208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1000_bdd_3_lut_23538.init = 16'hcaca;
    LUT4 n1000_bdd_3_lut_23697 (.A(n1000), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n31209)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1000_bdd_3_lut_23697.init = 16'he2e2;
    LUT4 Select_4184_i5_2_lut (.A(databus_out[10]), .B(rw), .Z(n5_adj_292)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4184_i5_2_lut.init = 16'h2222;
    LUT4 Select_4124_i5_2_lut (.A(databus_out[30]), .B(rw), .Z(n5_adj_300)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4124_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_346 (.A(\read_value[10]_adj_177 ), .B(read_value_adj_293[10]), 
         .C(n31716), .D(n46), .Z(n12_adj_295)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_346.init = 16'heca0;
    LUT4 i4_4_lut_adj_347 (.A(\read_value[30]_adj_178 ), .B(read_value_adj_293[30]), 
         .C(n31716), .D(n46), .Z(n12_adj_303)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_347.init = 16'heca0;
    LUT4 i7_4_lut_adj_348 (.A(n9_adj_309), .B(n14_adj_310), .C(n3_adj_179), 
         .D(n5_adj_312), .Z(databus[29])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_348.init = 16'hfffe;
    LUT4 register_addr_1__bdd_2_lut_23564 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n31228)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23564.init = 16'h2222;
    LUT4 i1_4_lut_adj_349 (.A(\read_value[29]_adj_180 ), .B(read_value[29]), 
         .C(n31719), .D(n47), .Z(n9_adj_309)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_349.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23565 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n31229)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23565.init = 16'he4e4;
    LUT4 i6_4_lut_adj_350 (.A(\read_value[29]_adj_181 ), .B(n12_adj_315), 
         .C(n6_adj_182), .D(n31703), .Z(n14_adj_310)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_350.init = 16'hfefc;
    LUT4 Select_4127_i5_2_lut (.A(databus_out[29]), .B(rw), .Z(n5_adj_312)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4127_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_351 (.A(\read_value[29]_adj_183 ), .B(read_value_adj_293[29]), 
         .C(n31716), .D(n46), .Z(n12_adj_315)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_351.init = 16'heca0;
    LUT4 i7_4_lut_adj_352 (.A(n9_adj_319), .B(n14_adj_320), .C(n3_adj_184), 
         .D(n5_adj_322), .Z(databus[9])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_352.init = 16'hfffe;
    LUT4 n1045_bdd_3_lut_23558 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n31231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1045_bdd_3_lut_23558.init = 16'hcaca;
    LUT4 i1_4_lut_adj_353 (.A(\read_value[9]_adj_185 ), .B(read_value[9]), 
         .C(n31719), .D(n47), .Z(n9_adj_319)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_353.init = 16'heca0;
    LUT4 i7_4_lut_adj_354 (.A(n9_adj_324), .B(n14_adj_325), .C(n3_adj_186), 
         .D(n5_adj_327), .Z(databus[28])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_354.init = 16'hfffe;
    LUT4 i1_4_lut_adj_355 (.A(\read_value[28]_adj_187 ), .B(read_value[28]), 
         .C(n31719), .D(n47), .Z(n9_adj_324)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_355.init = 16'heca0;
    LUT4 i6_4_lut_adj_356 (.A(\read_value[9]_adj_188 ), .B(n12_adj_330), 
         .C(n6_adj_189), .D(n31703), .Z(n14_adj_320)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_356.init = 16'hfefc;
    LUT4 n1045_bdd_3_lut_23659 (.A(n1045), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n31232)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1045_bdd_3_lut_23659.init = 16'he2e2;
    LUT4 i6_4_lut_adj_357 (.A(\read_value[28]_adj_190 ), .B(n12_adj_333), 
         .C(n6_adj_191), .D(n31703), .Z(n14_adj_325)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_357.init = 16'hfefc;
    LUT4 Select_4130_i5_2_lut (.A(databus_out[28]), .B(rw), .Z(n5_adj_327)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4130_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_358 (.A(\read_value[28]_adj_192 ), .B(read_value_adj_293[28]), 
         .C(n31716), .D(n46), .Z(n12_adj_333)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_358.init = 16'heca0;
    LUT4 Select_4187_i5_2_lut (.A(databus_out[9]), .B(rw), .Z(n5_adj_322)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4187_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_359 (.A(\read_value[9]_adj_193 ), .B(read_value_adj_293[9]), 
         .C(n31716), .D(n46), .Z(n12_adj_330)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_359.init = 16'heca0;
    LUT4 i7_4_lut_adj_360 (.A(n9_adj_339), .B(n14_adj_340), .C(n3_adj_194), 
         .D(n5_adj_342), .Z(databus[27])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_360.init = 16'hfffe;
    LUT4 i1_4_lut_adj_361 (.A(\read_value[27]_adj_195 ), .B(read_value[27]), 
         .C(n31719), .D(n47), .Z(n9_adj_339)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_361.init = 16'heca0;
    LUT4 i7_4_lut_adj_362 (.A(n9_adj_344), .B(n14_adj_345), .C(n3_adj_196), 
         .D(n5_adj_347), .Z(databus[8])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_362.init = 16'hfffe;
    LUT4 i6_4_lut_adj_363 (.A(\read_value[27]_adj_197 ), .B(n12_adj_349), 
         .C(n6_adj_198), .D(n31703), .Z(n14_adj_340)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_363.init = 16'hfefc;
    LUT4 Select_4133_i5_2_lut (.A(databus_out[27]), .B(n33446), .Z(n5_adj_342)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4133_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_364 (.A(\read_value[27]_adj_199 ), .B(read_value_adj_293[27]), 
         .C(n31716), .D(n46), .Z(n12_adj_349)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_364.init = 16'heca0;
    LUT4 i1_4_lut_adj_365 (.A(\read_value[8]_adj_200 ), .B(read_value[8]), 
         .C(n31719), .D(n47), .Z(n9_adj_344)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_365.init = 16'heca0;
    LUT4 i6_4_lut_adj_366 (.A(\read_value[8]_adj_201 ), .B(n12_adj_355), 
         .C(n6_adj_202), .D(n31703), .Z(n14_adj_345)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_366.init = 16'hfefc;
    LUT4 Select_4190_i5_2_lut (.A(databus_out[8]), .B(rw), .Z(n5_adj_347)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4190_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_367 (.A(\read_value[8]_adj_203 ), .B(read_value_adj_293[8]), 
         .C(n31716), .D(n46), .Z(n12_adj_355)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_367.init = 16'heca0;
    LUT4 i7_4_lut_adj_368 (.A(n9_adj_359), .B(n14_adj_360), .C(n3_adj_204), 
         .D(n5_adj_362), .Z(databus[26])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_368.init = 16'hfffe;
    LUT4 i1_4_lut_adj_369 (.A(\read_value[26]_adj_205 ), .B(read_value[26]), 
         .C(n31719), .D(n47), .Z(n9_adj_359)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_369.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23575 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n31243)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23575.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_23574 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n31242)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23574.init = 16'h2222;
    LUT4 i6_4_lut_adj_370 (.A(\read_value[26]_adj_206 ), .B(n12_adj_365), 
         .C(n6_adj_207), .D(n31703), .Z(n14_adj_360)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_370.init = 16'hfefc;
    LUT4 Select_4136_i5_2_lut (.A(databus_out[26]), .B(n33446), .Z(n5_adj_362)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4136_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_371 (.A(\read_value[26]_adj_208 ), .B(read_value_adj_293[26]), 
         .C(n31716), .D(n46), .Z(n12_adj_365)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_371.init = 16'heca0;
    PFUMX i23409 (.BLUT(n30838), .ALUT(n30837), .C0(\register_addr[1] ), 
          .Z(n30839));
    LUT4 i7_4_lut_adj_372 (.A(n9_adj_369), .B(n14_adj_370), .C(n3_adj_209), 
         .D(n5_adj_372), .Z(databus[25])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_372.init = 16'hfffe;
    LUT4 i1_4_lut_adj_373 (.A(\read_value[25]_adj_210 ), .B(read_value[25]), 
         .C(n31719), .D(n47), .Z(n9_adj_369)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_373.init = 16'heca0;
    LUT4 i6_4_lut_adj_374 (.A(\read_value[25]_adj_211 ), .B(n12_adj_375), 
         .C(n6_adj_212), .D(n31703), .Z(n14_adj_370)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_374.init = 16'hfefc;
    LUT4 \register_1[[5__bdd_3_lut_23644  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n31245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_23644 .init = 16'hcaca;
    LUT4 \register_1[[5__bdd_2_lut_23645  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n31246)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_23645 .init = 16'h8888;
    LUT4 Select_4139_i5_2_lut (.A(databus_out[25]), .B(n33446), .Z(n5_adj_372)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4139_i5_2_lut.init = 16'h2222;
    L6MUX21 i23357 (.D0(n30712), .D1(n30709), .SD(\register_addr[2] ), 
            .Z(n30713));
    LUT4 n1060_bdd_3_lut_23580 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n31271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1060_bdd_3_lut_23580.init = 16'hcaca;
    LUT4 n1060_bdd_3_lut_23629 (.A(n1060), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n31272)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1060_bdd_3_lut_23629.init = 16'he2e2;
    LUT4 i4_4_lut_adj_375 (.A(\read_value[25]_adj_213 ), .B(read_value_adj_293[25]), 
         .C(n31716), .D(n46), .Z(n12_adj_375)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_375.init = 16'heca0;
    LUT4 i1_4_lut_adj_376 (.A(\read_size[0] ), .B(\read_size[0]_adj_214 ), 
         .C(\select[2] ), .D(n31780), .Z(n9)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_376.init = 16'heca0;
    LUT4 i6_4_lut_adj_377 (.A(read_size_c[0]), .B(n12_adj_382), .C(n29694), 
         .D(\select[7] ), .Z(n14)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_377.init = 16'hfefc;
    LUT4 i7_4_lut_adj_378 (.A(n9_adj_384), .B(n14_adj_385), .C(n3_adj_215), 
         .D(n5_adj_387), .Z(databus[24])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_378.init = 16'hfffe;
    LUT4 i2_4_lut_adj_379 (.A(\select[4] ), .B(\read_size[0]_adj_216 ), 
         .C(n55), .D(n31762), .Z(n10)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_379.init = 16'heca0;
    LUT4 i4_4_lut_adj_380 (.A(read_size[0]), .B(n31732), .C(\select[1] ), 
         .D(\read_size[0]_adj_218 ), .Z(n12_adj_382)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_380.init = 16'heca0;
    LUT4 i5_4_lut (.A(n31741), .B(n10_adj_391), .C(n6_adj_219), .D(\read_size[2]_adj_220 ), 
         .Z(\reg_size[2] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfefc;
    LUT4 i4_4_lut_adj_381 (.A(n31732), .B(n8_adj_393), .C(n9_adj_221), 
         .D(\read_size[2]_adj_222 ), .Z(n10_adj_391)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_381.init = 16'hfefc;
    LUT4 i1_4_lut_adj_382 (.A(\read_value[24]_adj_223 ), .B(read_value[24]), 
         .C(n31719), .D(n47), .Z(n9_adj_384)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_382.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23678 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n31269)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23678.init = 16'he4e4;
    LUT4 i6_4_lut_adj_383 (.A(\read_value[24]_adj_224 ), .B(n12_adj_398), 
         .C(n6_adj_225), .D(n31703), .Z(n14_adj_385)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_383.init = 16'hfefc;
    LUT4 i2_4_lut_adj_384 (.A(read_size[2]), .B(\read_size[2]_adj_226 ), 
         .C(\select[1] ), .D(n31780), .Z(n8_adj_393)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_384.init = 16'heca0;
    LUT4 i9_4_lut (.A(n17), .B(n6_adj_402), .C(n16_adj_403), .D(n2), 
         .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 register_addr_1__bdd_2_lut_23677 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n31268)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23677.init = 16'h2222;
    LUT4 i7_4_lut_adj_385 (.A(\read_value[5]_adj_227 ), .B(n14_adj_404), 
         .C(n5), .D(n31719), .Z(n17)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_385.init = 16'hfefc;
    FD1S3IX read_value__i1 (.D(n31211), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n30843), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n31101), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n30713), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n31248), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(n31234), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i7 (.D(n31274), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 Select_4193_i6_2_lut (.A(databus_out[5]), .B(rw), .Z(n6_adj_402)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4193_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_386 (.A(read_value[5]), .B(n12_adj_408), .C(n8_adj_228), 
         .D(n47), .Z(n16_adj_403)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_386.init = 16'hfefc;
    LUT4 Select_4142_i5_2_lut (.A(databus_out[24]), .B(rw), .Z(n5_adj_387)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4142_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_387 (.A(\read_value[24]_adj_229 ), .B(read_value_adj_293[24]), 
         .C(n31716), .D(n46), .Z(n12_adj_398)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_387.init = 16'heca0;
    PFUMX i23355 (.BLUT(n30711), .ALUT(n30710), .C0(\register_addr[1] ), 
          .Z(n30712));
    LUT4 i7_4_lut_adj_388 (.A(n9_adj_412), .B(n14_adj_413), .C(n3_adj_230), 
         .D(n5_adj_415), .Z(databus[23])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_388.init = 16'hfffe;
    LUT4 i1_4_lut_adj_389 (.A(\read_value[23]_adj_231 ), .B(read_value[23]), 
         .C(n31719), .D(n47), .Z(n9_adj_412)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_389.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_23417 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n30838)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23417.init = 16'he4e4;
    LUT4 i6_4_lut_adj_390 (.A(\read_value[23]_adj_232 ), .B(n12_adj_418), 
         .C(n6_adj_233), .D(n31703), .Z(n14_adj_413)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_390.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_23416 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n30837)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23416.init = 16'h2222;
    LUT4 n1015_bdd_3_lut_23411 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n30840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1015_bdd_3_lut_23411.init = 16'hcaca;
    LUT4 Select_4145_i5_2_lut (.A(databus_out[23]), .B(n33446), .Z(n5_adj_415)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4145_i5_2_lut.init = 16'h2222;
    LUT4 i9_4_lut_adj_391 (.A(n17_adj_420), .B(n6_adj_421), .C(n16_adj_422), 
         .D(n2_adj_234), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_391.init = 16'hfffe;
    LUT4 i4_4_lut_adj_392 (.A(\read_value[23]_adj_235 ), .B(read_value_adj_293[23]), 
         .C(n31716), .D(n46), .Z(n12_adj_418)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_392.init = 16'heca0;
    LUT4 i4_4_lut_adj_393 (.A(read_value_adj_293[5]), .B(\read_value[5]_adj_236 ), 
         .C(n46), .D(n31733), .Z(n14_adj_404)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_393.init = 16'heca0;
    LUT4 i7_4_lut_adj_394 (.A(\read_value[6]_adj_237 ), .B(n14_adj_203), 
         .C(n5_adj_238), .D(n31719), .Z(n17_adj_420)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_394.init = 16'hfefc;
    LUT4 i7_4_lut_adj_395 (.A(n9_adj_430), .B(n14_adj_431), .C(n3_adj_239), 
         .D(n5_adj_433), .Z(databus[22])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_395.init = 16'hfffe;
    LUT4 i2_4_lut_adj_396 (.A(\read_value[5]_adj_240 ), .B(read_value_adj_538[5]), 
         .C(n31703), .D(n46_adj_208), .Z(n12_adj_408)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_396.init = 16'heca0;
    LUT4 i1_4_lut_adj_397 (.A(\read_value[22]_adj_241 ), .B(read_value[22]), 
         .C(n31719), .D(n47), .Z(n9_adj_430)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_397.init = 16'heca0;
    LUT4 i6_4_lut_adj_398 (.A(\read_value[22]_adj_242 ), .B(n12_adj_437), 
         .C(n6_adj_243), .D(n31703), .Z(n14_adj_431)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_398.init = 16'hfefc;
    LUT4 Select_4148_i5_2_lut (.A(databus_out[22]), .B(n33446), .Z(n5_adj_433)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4148_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_399 (.A(\read_value[22]_adj_244 ), .B(read_value_adj_293[22]), 
         .C(n31716), .D(n46), .Z(n12_adj_437)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_399.init = 16'heca0;
    LUT4 n1015_bdd_3_lut_23804 (.A(n1015), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n30841)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1015_bdd_3_lut_23804.init = 16'he2e2;
    LUT4 i7_4_lut_adj_400 (.A(n9_adj_441), .B(n14_adj_442), .C(n3_adj_245), 
         .D(n5_adj_444), .Z(databus[21])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_400.init = 16'hfffe;
    LUT4 i1_4_lut_adj_401 (.A(\read_value[21]_adj_246 ), .B(read_value[21]), 
         .C(n31719), .D(n47), .Z(n9_adj_441)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_401.init = 16'heca0;
    LUT4 i6_4_lut_adj_402 (.A(\read_value[21]_adj_247 ), .B(n12_adj_447), 
         .C(n6_adj_248), .D(n31703), .Z(n14_adj_442)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_402.init = 16'hfefc;
    LUT4 Select_4151_i5_2_lut (.A(databus_out[21]), .B(n33446), .Z(n5_adj_444)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4151_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_403 (.A(\read_value[21]_adj_249 ), .B(read_value_adj_293[21]), 
         .C(n31716), .D(n46), .Z(n12_adj_447)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_403.init = 16'heca0;
    LUT4 i7_4_lut_adj_404 (.A(n9_adj_451), .B(n14_adj_452), .C(n3_adj_250), 
         .D(n5_adj_454), .Z(databus[20])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_404.init = 16'hfffe;
    LUT4 Select_4207_i1_2_lut_rep_418 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n31841)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4207_i1_2_lut_rep_418.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n12795)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_4_lut_adj_405 (.A(\read_value[20]_adj_251 ), .B(read_value[20]), 
         .C(n31719), .D(n47), .Z(n9_adj_451)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_405.init = 16'heca0;
    LUT4 i6_4_lut_adj_406 (.A(\read_value[20]_adj_252 ), .B(n12_adj_457), 
         .C(n6_adj_253), .D(n31703), .Z(n14_adj_452)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_406.init = 16'hfefc;
    LUT4 Select_4192_i6_2_lut (.A(databus_out[6]), .B(rw), .Z(n6_adj_421)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4192_i6_2_lut.init = 16'h2222;
    LUT4 Select_4154_i5_2_lut (.A(databus_out[20]), .B(n33446), .Z(n5_adj_454)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4154_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_407 (.A(\read_value[20]_adj_254 ), .B(read_value_adj_293[20]), 
         .C(n31716), .D(n46), .Z(n12_adj_457)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_407.init = 16'heca0;
    L6MUX21 i23684 (.D0(n31562), .D1(n31559), .SD(\register_addr[2] ), 
            .Z(n31563));
    LUT4 i9_4_lut_adj_408 (.A(n17_adj_461), .B(n6_adj_462), .C(n16_adj_463), 
         .D(n2_adj_255), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_408.init = 16'hfffe;
    PFUMX i23682 (.BLUT(n31561), .ALUT(n31560), .C0(\register_addr[1] ), 
          .Z(n31562));
    LUT4 i7_4_lut_adj_409 (.A(n9_adj_465), .B(n14_adj_466), .C(n3_adj_256), 
         .D(n5_adj_468), .Z(databus[19])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_409.init = 16'hfffe;
    LUT4 i1_4_lut_adj_410 (.A(\read_value[19]_adj_257 ), .B(read_value[19]), 
         .C(n31719), .D(n47), .Z(n9_adj_465)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_410.init = 16'heca0;
    LUT4 i6_4_lut_adj_411 (.A(\read_value[19]_adj_258 ), .B(n12_adj_471), 
         .C(n6_adj_259), .D(n31703), .Z(n14_adj_466)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_411.init = 16'hfefc;
    LUT4 Select_4157_i5_2_lut (.A(databus_out[19]), .B(n33446), .Z(n5_adj_468)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4157_i5_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_412 (.A(\read_value[4]_adj_260 ), .B(n14_adj_474), 
         .C(n5_adj_261), .D(n31719), .Z(n17_adj_461)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_412.init = 16'hfefc;
    LUT4 i6_4_lut_adj_413 (.A(read_value[6]), .B(n12_adj_209), .C(n8_adj_262), 
         .D(n47), .Z(n16_adj_422)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_413.init = 16'hfefc;
    LUT4 Select_4194_i6_2_lut (.A(databus_out[4]), .B(n33446), .Z(n6_adj_462)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4194_i6_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_414 (.A(\read_value[19]_adj_263 ), .B(read_value_adj_293[19]), 
         .C(n31716), .D(n46), .Z(n12_adj_471)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_414.init = 16'heca0;
    PFUMX i23679 (.BLUT(n31558), .ALUT(n31557), .C0(\register_addr[1] ), 
          .Z(n31559));
    LUT4 i7_4_lut_adj_415 (.A(n9_c), .B(n14_c), .C(n3_adj_264), .D(n5_c), 
         .Z(databus[18])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_415.init = 16'hfffe;
    LUT4 i6_4_lut_adj_416 (.A(read_value[4]), .B(n12_adj_482), .C(n8_adj_265), 
         .D(n47), .Z(n16_adj_463)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_416.init = 16'hfefc;
    PFUMX i23353 (.BLUT(n30708), .ALUT(n30707), .C0(\register_addr[1] ), 
          .Z(n30709));
    LUT4 i4_4_lut_adj_417 (.A(read_value_adj_293[4]), .B(\read_value[4]_adj_266 ), 
         .C(n46), .D(n31733), .Z(n14_adj_474)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_417.init = 16'heca0;
    LUT4 i2_4_lut_adj_418 (.A(\read_value[4]_adj_267 ), .B(read_value_adj_538[4]), 
         .C(n31703), .D(n46_adj_208), .Z(n12_adj_482)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_418.init = 16'heca0;
    LUT4 i14_2_lut (.A(\select[7] ), .B(rw), .Z(n46_adj_208)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam i14_2_lut.init = 16'h8888;
    LUT4 i9_4_lut_adj_419 (.A(n17_adj_487), .B(n6_adj_488), .C(n16_adj_489), 
         .D(n2_adj_268), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_419.init = 16'hfffe;
    LUT4 i7_4_lut_adj_420 (.A(\read_value[3]_adj_269 ), .B(n14_adj_492), 
         .C(n5_adj_270), .D(n31719), .Z(n17_adj_487)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_420.init = 16'hfefc;
    LUT4 Select_4195_i6_2_lut (.A(databus_out[3]), .B(n33446), .Z(n6_adj_488)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4195_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_421 (.A(read_value[3]), .B(n12_adj_495), .C(n8_adj_271), 
         .D(n47), .Z(n16_adj_489)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_421.init = 16'hfefc;
    LUT4 i4_4_lut_adj_422 (.A(read_value_adj_293[3]), .B(\read_value[3]_adj_272 ), 
         .C(n46), .D(n31733), .Z(n14_adj_492)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_422.init = 16'heca0;
    FD1S3IX read_value__i0 (.D(n31563), .CK(\select[7] ), .CD(n31744), 
            .Q(read_value_adj_538[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=670, LSE_RLINE=682 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_423 (.A(\read_value[3]_adj_273 ), .B(read_value_adj_538[3]), 
         .C(n31703), .D(n46_adj_208), .Z(n12_adj_495)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_423.init = 16'heca0;
    LUT4 Select_4191_i6_2_lut (.A(databus_out[7]), .B(rw), .Z(n6_adj_501)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4191_i6_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_424 (.A(\read_value[7]_adj_274 ), .B(n14_adj_233), 
         .C(n5_adj_275), .D(n31719), .Z(n17_adj_504)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_424.init = 16'hfefc;
    LUT4 i1_4_lut_rep_321 (.A(\register_addr[2] ), .B(n29738), .C(\register_addr[0] ), 
         .D(\register_addr[1] ), .Z(n31744)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_rep_321.init = 16'heccc;
    L6MUX21 i23583 (.D0(n31273), .D1(n31270), .SD(\register_addr[2] ), 
            .Z(n31274));
    LUT4 i9_4_lut_adj_425 (.A(n17_adj_505), .B(n6_adj_506), .C(n16_adj_507), 
         .D(n2_adj_276), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_425.init = 16'hfffe;
    PFUMX i23578 (.BLUT(n31269), .ALUT(n31268), .C0(\register_addr[1] ), 
          .Z(n31270));
    PFUMX i23581 (.BLUT(n31272), .ALUT(n31271), .C0(\register_addr[1] ), 
          .Z(n31273));
    L6MUX21 i23572 (.D0(n31247), .D1(n31244), .SD(\register_addr[2] ), 
            .Z(n31248));
    PFUMX i23570 (.BLUT(n31246), .ALUT(n31245), .C0(\register_addr[1] ), 
          .Z(n31247));
    PFUMX i23568 (.BLUT(n31243), .ALUT(n31242), .C0(\register_addr[1] ), 
          .Z(n31244));
    LUT4 i7_4_lut_adj_426 (.A(\read_value[2]_adj_277 ), .B(n14_adj_510), 
         .C(n5_adj_278), .D(n31719), .Z(n17_adj_505)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_426.init = 16'hfefc;
    LUT4 i15547_1_lut_4_lut (.A(\register_addr[2] ), .B(n29738), .C(\register_addr[0] ), 
         .D(\register_addr[1] ), .Z(n176)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B))) */ ;
    defparam i15547_1_lut_4_lut.init = 16'h1333;
    LUT4 Select_4196_i6_2_lut (.A(databus_out[2]), .B(rw), .Z(n6_adj_506)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4196_i6_2_lut.init = 16'h2222;
    LUT4 i6_4_lut_adj_427 (.A(read_value[2]), .B(n12_adj_513), .C(n8_adj_279), 
         .D(n47), .Z(n16_adj_507)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_427.init = 16'hfefc;
    L6MUX21 i23561 (.D0(n31233), .D1(n31230), .SD(\register_addr[2] ), 
            .Z(n31234));
    PFUMX i23559 (.BLUT(n31232), .ALUT(n31231), .C0(\register_addr[1] ), 
          .Z(n31233));
    LUT4 i4_4_lut_adj_428 (.A(read_value_adj_293[2]), .B(\read_value[2]_adj_280 ), 
         .C(n46), .D(n31733), .Z(n14_adj_510)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_428.init = 16'heca0;
    PFUMX i23556 (.BLUT(n31229), .ALUT(n31228), .C0(\register_addr[1] ), 
          .Z(n31230));
    LUT4 i2_4_lut_adj_429 (.A(\read_value[2]_adj_281 ), .B(read_value_adj_538[2]), 
         .C(n31703), .D(n46_adj_208), .Z(n12_adj_513)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_429.init = 16'heca0;
    LUT4 i9_4_lut_adj_430 (.A(n1), .B(n18), .C(n14_adj_518), .D(n5_adj_282), 
         .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_430.init = 16'hfffe;
    L6MUX21 i23541 (.D0(n31210), .D1(n31207), .SD(\register_addr[2] ), 
            .Z(n31211));
    PFUMX i23539 (.BLUT(n31209), .ALUT(n31208), .C0(\register_addr[1] ), 
          .Z(n31210));
    PFUMX i23536 (.BLUT(n31206), .ALUT(n31205), .C0(\register_addr[1] ), 
          .Z(n31207));
    LUT4 i2_4_lut_adj_431 (.A(\read_value[0]_adj_283 ), .B(read_value_adj_538[0]), 
         .C(n31703), .D(n46_adj_208), .Z(n12_adj_242)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_431.init = 16'heca0;
    LUT4 i8_4_lut (.A(read_value_adj_293[1]), .B(n16_adj_522), .C(n2_adj_284), 
         .D(n46), .Z(n18)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut.init = 16'hfefc;
    LUT4 i4_4_lut_adj_432 (.A(read_value_adj_293[0]), .B(\read_value[0]_adj_285 ), 
         .C(n46), .D(n31733), .Z(n14_adj_526)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_432.init = 16'heca0;
    LUT4 i4_4_lut_adj_433 (.A(read_value[1]), .B(\read_value[1]_adj_286 ), 
         .C(n47), .D(n31733), .Z(n14_adj_518)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_433.init = 16'heca0;
    LUT4 i6_4_lut_adj_434 (.A(n11), .B(n4), .C(databus_out[1]), .D(n33446), 
         .Z(n16_adj_522)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i6_4_lut_adj_434.init = 16'heefe;
    LUT4 i9_4_lut_adj_435 (.A(n17_adj_504), .B(n6_adj_501), .C(n16), .D(n2_adj_287), 
         .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_435.init = 16'hfffe;
    LUT4 i1_4_lut_adj_436 (.A(\read_value[1]_adj_288 ), .B(read_value_adj_538[1]), 
         .C(n31746), .D(n46_adj_208), .Z(n11)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_436.init = 16'heca0;
    L6MUX21 i23499 (.D0(n31100), .D1(n31097), .SD(\register_addr[2] ), 
            .Z(n31101));
    PFUMX i23497 (.BLUT(n31099), .ALUT(n31098), .C0(\register_addr[1] ), 
          .Z(n31100));
    PFUMX i23494 (.BLUT(n31096), .ALUT(n31095), .C0(\register_addr[1] ), 
          .Z(n31097));
    LUT4 i9_4_lut_adj_437 (.A(n17_adj_531), .B(n6_adj_532), .C(n16_adj_244), 
         .D(n2_adj_289), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_437.init = 16'hfffe;
    LUT4 i7_4_lut_adj_438 (.A(\read_value[0]_adj_290 ), .B(n14_adj_526), 
         .C(n5_adj_291), .D(n31719), .Z(n17_adj_531)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_438.init = 16'hfefc;
    LUT4 Select_4198_i6_2_lut (.A(databus_out[0]), .B(n33446), .Z(n6_adj_532)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4198_i6_2_lut.init = 16'h2222;
    PWMReceiver recv_ch8 (.GND_net(GND_net), .debug_c_c(debug_c_c), .n31694(n31694), 
            .rc_ch8_c(rc_ch8_c), .n1060(n1060), .n27918(n27918), .n30160(n30160), 
            .n30216(n30216), .\register[6] ({\register[6] }), .n13719(n13719)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(257[14] 261[36])
    PWMReceiver_U1 recv_ch7 (.debug_c_c(debug_c_c), .n31694(n31694), .rc_ch7_c(rc_ch7_c), 
            .GND_net(GND_net), .n1045(n1045), .n27933(n27933), .n30195(n30195), 
            .\register[5] ({\register[5] }), .n14176(n14176), .n30205(n30205)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(252[14] 256[36])
    PWMReceiver_U2 recv_ch4 (.debug_c_c(debug_c_c), .n31694(n31694), .rc_ch4_c(rc_ch4_c), 
            .GND_net(GND_net), .n1030(n1030), .n27937(n27937), .n30182(n30182), 
            .\register[4] ({\register[4] }), .n14182(n14182), .n30191(n30191)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(247[14] 251[36])
    PWMReceiver_U3 recv_ch3 (.n30197(n30197), .debug_c_c(debug_c_c), .n31694(n31694), 
            .rc_ch3_c(rc_ch3_c), .GND_net(GND_net), .n1015(n1015), .n27924(n27924), 
            .\register[3] ({\register[3] }), .n14183(n14183), .n30189(n30189)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(242[14] 246[36])
    PWMReceiver_U4 recv_ch2 (.n30186(n30186), .GND_net(GND_net), .debug_c_c(debug_c_c), 
            .n31694(n31694), .rc_ch2_c(rc_ch2_c), .n1000(n1000), .n27915(n27915), 
            .\register[2] ({\register[2] }), .n14186(n14186), .n30218(n30218)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(237[14] 241[36])
    PWMReceiver_U5 recv_ch1 (.GND_net(GND_net), .debug_c_c(debug_c_c), .n31694(n31694), 
            .n29930(n29930), .\register[1] ({\register[1] }), .n14187(n14187), 
            .n9(n9_adj_292), .rc_ch1_c(rc_ch1_c), .n30152(n30152), .n30184(n30184), 
            .n985(n985), .n27912(n27912)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(232[17] 236[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (GND_net, debug_c_c, n31694, rc_ch8_c, n1060, n27918, 
            n30160, n30216, \register[6] , n13719) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n31694;
    input rc_ch8_c;
    output n1060;
    input n27918;
    output n30160;
    output n30216;
    output [7:0]\register[6] ;
    input n13719;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n31791;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31854, n31813, n29414, n31814, n29586, n28198, n1054, 
        n1066, n29906, n31857, n4, n28178, n26955, n31846;
    wire [15:0]n116;
    
    wire n26956, n31856, n28033, n6, n26954, n31855, n29990, n31858, 
        n31734, n26953, n13297, n31768, n29772, n28039, n33443, 
        n31767, n27230;
    wire [7:0]n958;
    
    wire n26958, n26957, n27229, n27228, n27227, n29587, n29691, 
        n10, n11, n16223;
    wire [7:0]n43;
    
    wire n26952, n27917, n5, n29947, n27952, n6_adj_190, n29773, 
        n26951;
    
    LUT4 i1_4_lut (.A(n31791), .B(count[8]), .C(n31854), .D(n31813), 
         .Z(n29414)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(count[4]), .B(n31814), .C(count[8]), .D(n29586), 
         .Z(n28198)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i22759_2_lut (.A(n1054), .B(n1066), .Z(n29906)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22759_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n31857), .D(n4), 
         .Z(n28178)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    CCU2D add_1740_11 (.A0(count[9]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31846), .C1(GND_net), .D1(GND_net), .CIN(n26955), 
          .COUT(n26956), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_11.INIT0 = 16'hd222;
    defparam add_1740_11.INIT1 = 16'hd222;
    defparam add_1740_11.INJECT1_0 = "NO";
    defparam add_1740_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_295 (.A(n31856), .B(count[9]), .C(n28033), .D(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_295.init = 16'heccc;
    LUT4 i2_4_lut_adj_296 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28033)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_296.init = 16'hfeee;
    CCU2D add_1740_9 (.A0(count[7]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31846), .C1(GND_net), .D1(GND_net), .CIN(n26954), 
          .COUT(n26955), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_9.INIT0 = 16'hd222;
    defparam add_1740_9.INIT1 = 16'hd222;
    defparam add_1740_9.INJECT1_0 = "NO";
    defparam add_1740_9.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_431 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n31854)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_431.init = 16'h8080;
    LUT4 i1_2_lut_rep_391_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n31814)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_391_4_lut.init = 16'h8000;
    LUT4 i15025_2_lut_rep_432 (.A(count[4]), .B(count[5]), .Z(n31855)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15025_2_lut_rep_432.init = 16'h8888;
    LUT4 i1_2_lut_rep_433 (.A(count[6]), .B(count[7]), .Z(n31856)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_433.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), .Z(n29586)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_rep_390_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[5]), 
         .D(count[4]), .Z(n31813)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_rep_390_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_434 (.A(count[11]), .B(count[10]), .Z(n31857)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_434.init = 16'heeee;
    LUT4 i22838_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n29990)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22838_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_435 (.A(count[15]), .B(count[14]), .Z(n31858)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_435.init = 16'heeee;
    LUT4 i1_2_lut_rep_311_3_lut (.A(count[15]), .B(count[14]), .C(n28178), 
         .Z(n31734)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_311_3_lut.init = 16'hfefe;
    CCU2D add_1740_7 (.A0(count[5]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31846), .C1(GND_net), .D1(GND_net), .CIN(n26953), 
          .COUT(n26954), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_7.INIT0 = 16'hd222;
    defparam add_1740_7.INIT1 = 16'hd222;
    defparam add_1740_7.INJECT1_0 = "NO";
    defparam add_1740_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_368 (.A(count[9]), .B(n13297), .Z(n31791)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_368.init = 16'heeee;
    LUT4 i1_2_lut_rep_345_3_lut (.A(count[9]), .B(n13297), .C(count[8]), 
         .Z(n31768)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_345_3_lut.init = 16'hfefe;
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n31694), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1066));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1066), .SP(n31694), .CK(debug_c_c), .Q(n1054));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    FD1P3AX valid_48 (.D(n29772), .SP(n27918), .CK(debug_c_c), .Q(n1060));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i15626_3_lut_rep_450 (.A(n28039), .B(n13297), .C(count[9]), .Z(n33443)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15626_3_lut_rep_450.init = 16'hecec;
    LUT4 i21_3_lut_rep_344_4_lut_4_lut (.A(n28039), .B(n13297), .C(count[9]), 
         .D(n28198), .Z(n31767)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i21_3_lut_rep_344_4_lut_4_lut.init = 16'h1310;
    CCU2D sub_65_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27230), 
          .S0(n958[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_9.INIT1 = 16'h0000;
    defparam sub_65_add_2_9.INJECT1_0 = "NO";
    defparam sub_65_add_2_9.INJECT1_1 = "NO";
    CCU2D add_1740_17 (.A0(count[15]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26958), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_17.INIT0 = 16'hd222;
    defparam add_1740_17.INIT1 = 16'h0000;
    defparam add_1740_17.INJECT1_0 = "NO";
    defparam add_1740_17.INJECT1_1 = "NO";
    CCU2D add_1740_15 (.A0(count[13]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31846), .C1(GND_net), .D1(GND_net), .CIN(n26957), 
          .COUT(n26958), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_15.INIT0 = 16'hd222;
    defparam add_1740_15.INIT1 = 16'hd222;
    defparam add_1740_15.INJECT1_0 = "NO";
    defparam add_1740_15.INJECT1_1 = "NO";
    CCU2D sub_65_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27229), 
          .COUT(n27230), .S0(n958[5]), .S1(n958[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_65_add_2_7.INJECT1_0 = "NO";
    defparam sub_65_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_65_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27228), 
          .COUT(n27229), .S0(n958[3]), .S1(n958[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_65_add_2_5.INJECT1_0 = "NO";
    defparam sub_65_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_65_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27227), 
          .COUT(n27228), .S0(n958[1]), .S1(n958[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_65_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_65_add_2_3.INJECT1_0 = "NO";
    defparam sub_65_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_65_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27227), 
          .S1(n958[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_65_add_2_1.INIT0 = 16'hF000;
    defparam sub_65_add_2_1.INIT1 = 16'h5555;
    defparam sub_65_add_2_1.INJECT1_0 = "NO";
    defparam sub_65_add_2_1.INJECT1_1 = "NO";
    LUT4 i23209_3_lut_3_lut_4_lut (.A(n29587), .B(n31768), .C(n33443), 
         .D(n31734), .Z(n29772)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23209_3_lut_3_lut_4_lut.init = 16'h000e;
    CCU2D add_1740_13 (.A0(count[11]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31846), .C1(GND_net), .D1(GND_net), .CIN(n26956), 
          .COUT(n26957), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_13.INIT0 = 16'hd222;
    defparam add_1740_13.INIT1 = 16'hd222;
    defparam add_1740_13.INJECT1_0 = "NO";
    defparam add_1740_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[0]), .B(n31854), .C(n31856), .D(n31855), 
         .Z(n29691)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23105_4_lut (.A(n31767), .B(n29906), .C(n29414), .D(n10), 
         .Z(n30160)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23105_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_297 (.A(n31694), .B(n31858), .C(n11), .D(n29990), 
         .Z(n16223)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_297.init = 16'h0020;
    LUT4 i4_4_lut (.A(n28198), .B(n29906), .C(n28039), .D(count[9]), 
         .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i15102_2_lut (.A(n958[0]), .B(n29414), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15102_2_lut.init = 16'h2222;
    CCU2D add_1740_5 (.A0(count[3]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31846), .C1(GND_net), .D1(GND_net), .CIN(n26952), 
          .COUT(n26953), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_5.INIT0 = 16'hd222;
    defparam add_1740_5.INIT1 = 16'hd222;
    defparam add_1740_5.INJECT1_0 = "NO";
    defparam add_1740_5.INJECT1_1 = "NO";
    LUT4 i15343_2_lut (.A(n958[7]), .B(n29414), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15343_2_lut.init = 16'h2222;
    LUT4 i15342_2_lut (.A(n958[6]), .B(n29414), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15342_2_lut.init = 16'h2222;
    LUT4 i15341_2_lut (.A(n958[5]), .B(n29414), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15341_2_lut.init = 16'h2222;
    LUT4 i15340_2_lut (.A(n958[4]), .B(n29414), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15340_2_lut.init = 16'h2222;
    LUT4 i15339_2_lut (.A(n958[3]), .B(n29414), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15339_2_lut.init = 16'h2222;
    LUT4 i15338_2_lut (.A(n958[2]), .B(n29414), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15338_2_lut.init = 16'h2222;
    LUT4 i15337_2_lut (.A(n958[1]), .B(n29414), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15337_2_lut.init = 16'h2222;
    LUT4 i23161_4_lut (.A(n31858), .B(n31846), .C(n28178), .D(n27917), 
         .Z(n30216)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23161_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_298 (.A(n5), .B(n29906), .C(n29947), .D(n33443), 
         .Z(n27917)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_298.init = 16'hccec;
    LUT4 i3_4_lut_adj_299 (.A(n27952), .B(n6_adj_190), .C(count[8]), .D(n31855), 
         .Z(n28039)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_299.init = 16'hfefc;
    LUT4 i3_4_lut_adj_300 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27952)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_300.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6_adj_190)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_301 (.A(count[12]), .B(count[13]), .C(n31858), .D(n31857), 
         .Z(n13297)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_301.init = 16'hfffe;
    LUT4 i1_4_lut_adj_302 (.A(count[4]), .B(n29586), .C(count[3]), .D(n6), 
         .Z(n29587)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_302.init = 16'hccc8;
    LUT4 i2899_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2899_2_lut.init = 16'h8888;
    LUT4 i5_2_lut_rep_423 (.A(n1054), .B(n1066), .Z(n31846)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_423.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_303 (.A(n1054), .B(n1066), .C(n28178), 
         .D(n31858), .Z(n29773)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_4_lut_adj_303.init = 16'hfff4;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13719), .PD(n16223), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1740_3 (.A0(count[1]), .B0(n31846), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31846), .C1(GND_net), .D1(GND_net), .CIN(n26951), 
          .COUT(n26952), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_3.INIT0 = 16'hd222;
    defparam add_1740_3.INIT1 = 16'hd222;
    defparam add_1740_3.INJECT1_0 = "NO";
    defparam add_1740_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(n28198), .B(n33443), .C(n31791), .D(n29414), 
         .Z(n5)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    LUT4 i22795_3_lut_4_lut (.A(count[8]), .B(n31791), .C(n29587), .D(n29691), 
         .Z(n29947)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22795_3_lut_4_lut.init = 16'hfeee;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31791), .C(n29691), 
         .D(n29587), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    CCU2D add_1740_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29773), .B1(n1066), .C1(count[0]), .D1(n1054), .COUT(n26951), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1740_1.INIT0 = 16'hF000;
    defparam add_1740_1.INIT1 = 16'ha565;
    defparam add_1740_1.INJECT1_0 = "NO";
    defparam add_1740_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (debug_c_c, n31694, rc_ch7_c, GND_net, n1045, 
            n27933, n30195, \register[5] , n14176, n30205) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31694;
    input rc_ch7_c;
    input GND_net;
    output n1045;
    input n27933;
    output n30195;
    output [7:0]\register[5] ;
    input n14176;
    output n30205;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n29598, n31764, n33441, n31735, n29719;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31849, n29389, n31850, n31810, n31859, n30002, n31860, 
        n29597, n31861, n28179, n5, n29718, n29412;
    wire [7:0]n949;
    wire [7:0]n43;
    
    wire n28043, n13338, n31788, n1051, n1039, n26961;
    wire [15:0]n116;
    
    wire n26962, n26960, n26959, n28199, n31761, n27234, n27233, 
        n27232, n27231, n27930, n5_adj_188, n29729, n29941, n6, 
        n29669, n26966, n26965, n27899, n6_adj_189, n26964, n26963, 
        n16117, n4, n28087, n10, n11, n8;
    
    LUT4 i23211_3_lut_3_lut_4_lut (.A(n29598), .B(n31764), .C(n33441), 
         .D(n31735), .Z(n29719)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23211_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i2_3_lut_rep_426 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n31849)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_rep_426.init = 16'h8080;
    LUT4 i1_2_lut_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), .D(count[0]), 
         .Z(n29389)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i14644_2_lut_rep_427 (.A(count[4]), .B(count[5]), .Z(n31850)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14644_2_lut_rep_427.init = 16'h8888;
    LUT4 i2_3_lut_rep_387_4_lut (.A(count[4]), .B(count[5]), .C(count[7]), 
         .D(count[6]), .Z(n31810)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_387_4_lut.init = 16'h8000;
    LUT4 i22747_2_lut_rep_436 (.A(count[11]), .B(count[10]), .Z(n31859)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22747_2_lut_rep_436.init = 16'heeee;
    LUT4 i22850_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n30002)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22850_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_437 (.A(count[6]), .B(count[7]), .Z(n31860)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_437.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), .Z(n29597)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_438 (.A(count[15]), .B(count[14]), .Z(n31861)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_438.init = 16'heeee;
    LUT4 i1_2_lut_rep_312_3_lut (.A(count[15]), .B(count[14]), .C(n28179), 
         .Z(n31735)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_312_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n28179), 
         .Z(n29718)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(n29412), .B(n949[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_adj_276 (.A(n29412), .B(n949[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_276.init = 16'h4444;
    LUT4 i15590_3_lut_rep_448 (.A(n28043), .B(n13338), .C(count[9]), .Z(n33441)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15590_3_lut_rep_448.init = 16'hecec;
    LUT4 i1_2_lut_rep_365 (.A(count[9]), .B(n13338), .Z(n31788)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_365.init = 16'heeee;
    LUT4 i1_2_lut_rep_341_3_lut (.A(count[9]), .B(n13338), .C(count[8]), 
         .Z(n31764)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_341_3_lut.init = 16'hfefe;
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n31694), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1051));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1051), .SP(n31694), .CK(debug_c_c), .Q(n1039));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D add_1736_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26961), 
          .COUT(n26962), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_7.INIT0 = 16'hd222;
    defparam add_1736_7.INIT1 = 16'hd222;
    defparam add_1736_7.INJECT1_0 = "NO";
    defparam add_1736_7.INJECT1_1 = "NO";
    CCU2D add_1736_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26960), 
          .COUT(n26961), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_5.INIT0 = 16'hd222;
    defparam add_1736_5.INIT1 = 16'hd222;
    defparam add_1736_5.INJECT1_0 = "NO";
    defparam add_1736_5.INJECT1_1 = "NO";
    CCU2D add_1736_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26959), 
          .COUT(n26960), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_3.INIT0 = 16'hd222;
    defparam add_1736_3.INIT1 = 16'hd222;
    defparam add_1736_3.INJECT1_0 = "NO";
    defparam add_1736_3.INJECT1_1 = "NO";
    LUT4 i21_3_lut_rep_338_4_lut_4_lut (.A(n28043), .B(n13338), .C(count[9]), 
         .D(n28199), .Z(n31761)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i21_3_lut_rep_338_4_lut_4_lut.init = 16'h1310;
    CCU2D add_1736_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29718), .B1(n1051), .C1(count[0]), .D1(n1039), .COUT(n26959), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_1.INIT0 = 16'hF000;
    defparam add_1736_1.INIT1 = 16'ha565;
    defparam add_1736_1.INJECT1_0 = "NO";
    defparam add_1736_1.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27234), 
          .S0(n949[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_9.INIT1 = 16'h0000;
    defparam sub_64_add_2_9.INJECT1_0 = "NO";
    defparam sub_64_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27233), 
          .COUT(n27234), .S0(n949[5]), .S1(n949[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_64_add_2_7.INJECT1_0 = "NO";
    defparam sub_64_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27232), 
          .COUT(n27233), .S0(n949[3]), .S1(n949[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_64_add_2_5.INJECT1_0 = "NO";
    defparam sub_64_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27231), 
          .COUT(n27232), .S0(n949[1]), .S1(n949[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_64_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_64_add_2_3.INJECT1_0 = "NO";
    defparam sub_64_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_64_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27231), 
          .S1(n949[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_64_add_2_1.INIT0 = 16'hF000;
    defparam sub_64_add_2_1.INIT1 = 16'h5555;
    defparam sub_64_add_2_1.INJECT1_0 = "NO";
    defparam sub_64_add_2_1.INJECT1_1 = "NO";
    FD1P3AX valid_48 (.D(n29719), .SP(n27933), .CK(debug_c_c), .Q(n1045));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i23140_4_lut (.A(n31861), .B(n5), .C(n28179), .D(n27930), .Z(n30195)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23140_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5_adj_188), .B(n29729), .C(n29941), .D(n33441), 
         .Z(n27930)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i1_4_lut_adj_277 (.A(count[4]), .B(n29597), .C(count[3]), .D(n6), 
         .Z(n29598)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_277.init = 16'hccc8;
    LUT4 i1_2_lut_4_lut_adj_278 (.A(count[6]), .B(count[7]), .C(n31850), 
         .D(n29389), .Z(n29669)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_278.init = 16'h8000;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n31861), .D(n31859), 
         .Z(n13338)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_279 (.A(n31788), .B(count[8]), .C(n31849), .D(n31810), 
         .Z(n29412)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_279.init = 16'hfbbb;
    CCU2D add_1736_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26966), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_17.INIT0 = 16'hd222;
    defparam add_1736_17.INIT1 = 16'h0000;
    defparam add_1736_17.INJECT1_0 = "NO";
    defparam add_1736_17.INJECT1_1 = "NO";
    CCU2D add_1736_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26965), 
          .COUT(n26966), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_15.INIT0 = 16'hd222;
    defparam add_1736_15.INIT1 = 16'hd222;
    defparam add_1736_15.INJECT1_0 = "NO";
    defparam add_1736_15.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_280 (.A(count[4]), .B(n29389), .C(count[8]), .D(n29597), 
         .Z(n28199)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_280.init = 16'h8000;
    LUT4 i1_2_lut_adj_281 (.A(n1051), .B(n1039), .Z(n29729)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_281.init = 16'hbbbb;
    LUT4 i3_4_lut_adj_282 (.A(n27899), .B(n6_adj_189), .C(count[8]), .D(n31850), 
         .Z(n28043)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_282.init = 16'hfefc;
    LUT4 i3_4_lut_adj_283 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27899)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_283.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6_adj_189)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i5_2_lut (.A(n1039), .B(n1051), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    CCU2D add_1736_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26964), 
          .COUT(n26965), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_13.INIT0 = 16'hd222;
    defparam add_1736_13.INIT1 = 16'hd222;
    defparam add_1736_13.INJECT1_0 = "NO";
    defparam add_1736_13.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    CCU2D add_1736_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26963), 
          .COUT(n26964), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_11.INIT0 = 16'hd222;
    defparam add_1736_11.INIT1 = 16'hd222;
    defparam add_1736_11.INJECT1_0 = "NO";
    defparam add_1736_11.INJECT1_1 = "NO";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    CCU2D add_1736_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26962), 
          .COUT(n26963), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1736_9.INIT0 = 16'hd222;
    defparam add_1736_9.INIT1 = 16'hd222;
    defparam add_1736_9.INJECT1_0 = "NO";
    defparam add_1736_9.INJECT1_1 = "NO";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n31859), .D(n4), 
         .Z(n28179)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_284 (.A(n31860), .B(count[9]), .C(n28087), .D(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_284.init = 16'heccc;
    LUT4 i2_4_lut_adj_285 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28087)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_285.init = 16'hfeee;
    LUT4 i2957_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2957_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_286 (.A(n29412), .B(n949[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_286.init = 16'h4444;
    LUT4 i1_2_lut_adj_287 (.A(n29412), .B(n949[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_287.init = 16'h4444;
    LUT4 i1_2_lut_adj_288 (.A(n29412), .B(n949[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_288.init = 16'h4444;
    LUT4 i1_2_lut_adj_289 (.A(n29412), .B(n949[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_289.init = 16'h4444;
    LUT4 i1_2_lut_4_lut_adj_290 (.A(n28199), .B(n33441), .C(n31788), .D(n29412), 
         .Z(n5_adj_188)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut_adj_290.init = 16'hcd00;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31788), .C(n29669), 
         .D(n29598), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22791_3_lut_4_lut (.A(count[8]), .B(n31788), .C(n29598), .D(n29669), 
         .Z(n29941)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i22791_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_adj_291 (.A(n29412), .B(n949[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_291.init = 16'h4444;
    LUT4 i1_2_lut_adj_292 (.A(n29412), .B(n949[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_292.init = 16'h4444;
    LUT4 i23150_4_lut (.A(n31761), .B(n29729), .C(n29412), .D(n10), 
         .Z(n30205)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23150_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_293 (.A(n31694), .B(n31861), .C(n11), .D(n30002), 
         .Z(n16117)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_293.init = 16'h0020;
    LUT4 i4_4_lut (.A(n28199), .B(n8), .C(n28043), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0c88;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14176), .PD(n16117), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_294 (.A(n1039), .B(n1051), .Z(n8)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_adj_294.init = 16'h2222;
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (debug_c_c, n31694, rc_ch4_c, GND_net, n1030, 
            n27937, n30182, \register[4] , n14182, n30191) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31694;
    input rc_ch4_c;
    input GND_net;
    output n1030;
    input n27937;
    output n30182;
    output [7:0]\register[4] ;
    input n14182;
    output n30191;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n4, n4_adj_184, n31847, n31809, n13367, n28037, n10, 
        n31758, n1024, n1036, n31786, n31760, n26974, n5;
    wire [15:0]n116;
    
    wire n26973, n27238;
    wire [7:0]n940;
    
    wire n27237, n27236, n27235, n26972, n26971, n26970, n26969, 
        n29748, n31845, n29395, n29601, n26968, n26967, n29749, 
        n31844, n28180, n27936, n33440, n29898, n7, n29822, n31843, 
        n27901, n6, n27774, n16122;
    wire [7:0]n43;
    
    wire n31842, n4_adj_185, n4_adj_186, n31808, n30000, n31729, 
        n10_adj_187, n11;
    
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_184)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i14769_2_lut_rep_424 (.A(count[4]), .B(count[5]), .Z(n31847)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14769_2_lut_rep_424.init = 16'h8888;
    LUT4 i2_3_lut_rep_386_4_lut (.A(count[4]), .B(count[5]), .C(count[6]), 
         .D(count[7]), .Z(n31809)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_386_4_lut.init = 16'h8000;
    LUT4 i21_3_lut_rep_335_4_lut_4_lut (.A(n13367), .B(n28037), .C(count[9]), 
         .D(n10), .Z(n31758)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam i21_3_lut_rep_335_4_lut_4_lut.init = 16'h1510;
    FD1P3AX prev_in_46 (.D(n1036), .SP(n31694), .CK(debug_c_c), .Q(n1024));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_363 (.A(count[9]), .B(n13367), .Z(n31786)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_363.init = 16'heeee;
    LUT4 i1_2_lut_rep_337_3_lut (.A(count[9]), .B(n13367), .C(count[8]), 
         .Z(n31760)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_337_3_lut.init = 16'hfefe;
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n31694), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1036));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    CCU2D add_1732_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26974), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_17.INIT0 = 16'hd222;
    defparam add_1732_17.INIT1 = 16'h0000;
    defparam add_1732_17.INJECT1_0 = "NO";
    defparam add_1732_17.INJECT1_1 = "NO";
    CCU2D add_1732_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26973), 
          .COUT(n26974), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_15.INIT0 = 16'hd222;
    defparam add_1732_15.INIT1 = 16'hd222;
    defparam add_1732_15.INJECT1_0 = "NO";
    defparam add_1732_15.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27238), 
          .S0(n940[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_9.INIT1 = 16'h0000;
    defparam sub_63_add_2_9.INJECT1_0 = "NO";
    defparam sub_63_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27237), 
          .COUT(n27238), .S0(n940[5]), .S1(n940[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_63_add_2_7.INJECT1_0 = "NO";
    defparam sub_63_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27236), 
          .COUT(n27237), .S0(n940[3]), .S1(n940[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_63_add_2_5.INJECT1_0 = "NO";
    defparam sub_63_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27235), 
          .COUT(n27236), .S0(n940[1]), .S1(n940[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_63_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_63_add_2_3.INJECT1_0 = "NO";
    defparam sub_63_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_63_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27235), 
          .S1(n940[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_63_add_2_1.INIT0 = 16'hF000;
    defparam sub_63_add_2_1.INIT1 = 16'h5555;
    defparam sub_63_add_2_1.INJECT1_0 = "NO";
    defparam sub_63_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1732_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26972), 
          .COUT(n26973), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_13.INIT0 = 16'hd222;
    defparam add_1732_13.INIT1 = 16'hd222;
    defparam add_1732_13.INJECT1_0 = "NO";
    defparam add_1732_13.INJECT1_1 = "NO";
    CCU2D add_1732_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26971), 
          .COUT(n26972), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_11.INIT0 = 16'hd222;
    defparam add_1732_11.INIT1 = 16'hd222;
    defparam add_1732_11.INJECT1_0 = "NO";
    defparam add_1732_11.INJECT1_1 = "NO";
    CCU2D add_1732_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26970), 
          .COUT(n26971), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_9.INIT0 = 16'hd222;
    defparam add_1732_9.INIT1 = 16'hd222;
    defparam add_1732_9.INJECT1_0 = "NO";
    defparam add_1732_9.INJECT1_1 = "NO";
    CCU2D add_1732_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26969), 
          .COUT(n26970), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_7.INIT0 = 16'hd222;
    defparam add_1732_7.INIT1 = 16'hd222;
    defparam add_1732_7.INJECT1_0 = "NO";
    defparam add_1732_7.INJECT1_1 = "NO";
    FD1P3AX valid_48 (.D(n29748), .SP(n27937), .CK(debug_c_c), .Q(n1030));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i3_3_lut_4_lut (.A(count[8]), .B(n31845), .C(n29395), .D(n31847), 
         .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut (.A(count[7]), .B(count[6]), .C(n31847), .D(n29395), 
         .Z(n29601)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8000;
    CCU2D add_1732_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26968), 
          .COUT(n26969), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_5.INIT0 = 16'hd222;
    defparam add_1732_5.INIT1 = 16'hd222;
    defparam add_1732_5.INJECT1_0 = "NO";
    defparam add_1732_5.INJECT1_1 = "NO";
    CCU2D add_1732_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26967), 
          .COUT(n26968), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_3.INIT0 = 16'hd222;
    defparam add_1732_3.INIT1 = 16'hd222;
    defparam add_1732_3.INJECT1_0 = "NO";
    defparam add_1732_3.INJECT1_1 = "NO";
    CCU2D add_1732_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29749), .B1(n1036), .C1(count[0]), .D1(n1024), .COUT(n26967), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1732_1.INIT0 = 16'hF000;
    defparam add_1732_1.INIT1 = 16'ha565;
    defparam add_1732_1.INJECT1_0 = "NO";
    defparam add_1732_1.INJECT1_1 = "NO";
    LUT4 i23127_4_lut (.A(n31844), .B(n5), .C(n28180), .D(n27936), .Z(n30182)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23127_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n33440), .B(n29898), .C(n7), .D(n29822), .Z(n27936)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n31844), .D(n31843), 
         .Z(n13367)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_261 (.A(n27901), .B(n6), .C(count[8]), .D(n31847), 
         .Z(n28037)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_261.init = 16'hfefc;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_262 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27901)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_262.init = 16'hfffe;
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(n31845), .B(count[4]), .C(count[5]), .D(n4), .Z(n27774)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_263 (.A(n31809), .B(n31786), .C(n31842), .D(count[8]), 
         .Z(n4_adj_185)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_263.init = 16'hecff;
    LUT4 i22751_2_lut (.A(n1024), .B(n1036), .Z(n29898)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22751_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_adj_264 (.A(count[13]), .B(count[12]), .C(n31843), .D(n4_adj_186), 
         .Z(n28180)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_264.init = 16'h8880;
    LUT4 i1_4_lut_adj_265 (.A(count[9]), .B(count[5]), .C(n31808), .D(n4_adj_184), 
         .Z(n4_adj_186)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_265.init = 16'hfaea;
    LUT4 i22675_3_lut_rep_447 (.A(n13367), .B(n28037), .C(count[9]), .Z(n33440)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i22675_3_lut_rep_447.init = 16'heaea;
    LUT4 i5_2_lut (.A(n1024), .B(n1036), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_rep_419 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n31842)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_rep_419.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_266 (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n29395)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_4_lut_adj_266.init = 16'h8000;
    LUT4 i22743_2_lut_rep_420 (.A(count[11]), .B(count[10]), .Z(n31843)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22743_2_lut_rep_420.init = 16'heeee;
    LUT4 i22848_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n30000)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22848_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_421 (.A(count[15]), .B(count[14]), .Z(n31844)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_421.init = 16'heeee;
    LUT4 i1_2_lut_rep_306_3_lut (.A(count[15]), .B(count[14]), .C(n28180), 
         .Z(n31729)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_306_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n28180), 
         .Z(n29749)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_422 (.A(count[6]), .B(count[7]), .Z(n31845)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_422.init = 16'h8888;
    LUT4 i23207_3_lut_3_lut_4_lut (.A(n27774), .B(n31760), .C(n33440), 
         .D(n31729), .Z(n29748)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23207_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_2_lut_rep_385_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n31808)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_385_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(n4_adj_185), .B(n940[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_4_lut_adj_267 (.A(n10), .B(n33440), .C(n31786), .D(n4_adj_185), 
         .Z(n7)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut_adj_267.init = 16'hcd00;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31786), .C(n29601), 
         .D(n27774), .Z(n10_adj_187)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22677_3_lut_4_lut (.A(count[8]), .B(n31786), .C(n27774), .D(n29601), 
         .Z(n29822)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22677_3_lut_4_lut.init = 16'hfeee;
    LUT4 i23136_4_lut (.A(n31758), .B(n29898), .C(n4_adj_185), .D(n10_adj_187), 
         .Z(n30191)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23136_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_268 (.A(n31694), .B(n31844), .C(n11), .D(n30000), 
         .Z(n16122)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_268.init = 16'h0020;
    LUT4 i4_4_lut (.A(n10), .B(n29898), .C(n28037), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i1_2_lut_adj_269 (.A(n4_adj_185), .B(n940[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_269.init = 16'h4444;
    LUT4 i1_2_lut_adj_270 (.A(n4_adj_185), .B(n940[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_270.init = 16'h4444;
    LUT4 i1_2_lut_adj_271 (.A(n4_adj_185), .B(n940[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_271.init = 16'h4444;
    LUT4 i1_2_lut_adj_272 (.A(n4_adj_185), .B(n940[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_272.init = 16'h4444;
    LUT4 i1_2_lut_adj_273 (.A(n4_adj_185), .B(n940[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_273.init = 16'h4444;
    LUT4 i1_2_lut_adj_274 (.A(n4_adj_185), .B(n940[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_274.init = 16'h4444;
    LUT4 i1_2_lut_adj_275 (.A(n4_adj_185), .B(n940[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_275.init = 16'h4444;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14182), .PD(n16122), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (n30197, debug_c_c, n31694, rc_ch3_c, GND_net, 
            n1015, n27924, \register[3] , n14183, n30189) /* synthesis syn_module_defined=1 */ ;
    output n30197;
    input debug_c_c;
    input n31694;
    input rc_ch3_c;
    input GND_net;
    output n1015;
    input n27924;
    output [7:0]\register[3] ;
    input n14183;
    output n30189;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n28201, n33442, n31766, n29416, n5;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31851, n29381, n31852, n31811, n29697, n29512, n10, 
        n29945, n31868, n29511, n31869, n28181, n31740, n31812, 
        n5_adj_182, n29779, n29759, n27923, n29864, n1021, n26975;
    wire [15:0]n116;
    
    wire n26976, n1009, n27242;
    wire [7:0]n931;
    
    wire n27241, n27240, n27239, n27970, n31789, n31731, n29778, 
        n6, n31730, n28061, n6_adj_183, n4, n28007, n26982, n16124;
    wire [7:0]n43;
    
    wire n26981, n26980, n26979, n26978, n26977, n16, n26;
    
    LUT4 i1_2_lut_4_lut (.A(n28201), .B(n33442), .C(n31766), .D(n29416), 
         .Z(n5)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    LUT4 i2_3_lut_rep_428 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n31851)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_rep_428.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_245 (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n29381)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_4_lut_adj_245.init = 16'h8000;
    LUT4 i15297_2_lut_rep_429 (.A(count[4]), .B(count[5]), .Z(n31852)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15297_2_lut_rep_429.init = 16'h8888;
    LUT4 i2_3_lut_rep_388_4_lut (.A(count[4]), .B(count[5]), .C(count[6]), 
         .D(count[7]), .Z(n31811)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_388_4_lut.init = 16'h8000;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31766), .C(n29697), 
         .D(n29512), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22794_3_lut_4_lut (.A(count[8]), .B(n31766), .C(n29512), .D(n29697), 
         .Z(n29945)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22794_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_rep_445 (.A(count[6]), .B(count[7]), .Z(n31868)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_445.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), .Z(n29511)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_446 (.A(count[15]), .B(count[14]), .Z(n31869)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_446.init = 16'heeee;
    LUT4 i1_2_lut_rep_317_3_lut (.A(count[15]), .B(count[14]), .C(n28181), 
         .Z(n31740)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_317_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_389_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n31812)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_389_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5_adj_182), 
         .D(n28181), .Z(n29779)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_343_4_lut (.A(n31812), .B(count[13]), .C(n29759), 
         .D(count[9]), .Z(n31766)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_343_4_lut.init = 16'hfffe;
    LUT4 i23142_4_lut (.A(n31869), .B(n5_adj_182), .C(n28181), .D(n27923), 
         .Z(n30197)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23142_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5), .B(n29864), .C(n29945), .D(n33442), .Z(n27923)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n31694), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1021));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    CCU2D add_1728_3 (.A0(count[1]), .B0(n5_adj_182), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5_adj_182), .C1(GND_net), .D1(GND_net), 
          .CIN(n26975), .COUT(n26976), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_3.INIT0 = 16'hd222;
    defparam add_1728_3.INIT1 = 16'hd222;
    defparam add_1728_3.INJECT1_0 = "NO";
    defparam add_1728_3.INJECT1_1 = "NO";
    CCU2D add_1728_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29779), .B1(n1021), .C1(count[0]), .D1(n1009), .COUT(n26975), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_1.INIT0 = 16'hF000;
    defparam add_1728_1.INIT1 = 16'ha565;
    defparam add_1728_1.INJECT1_0 = "NO";
    defparam add_1728_1.INJECT1_1 = "NO";
    FD1P3AX prev_in_46 (.D(n1021), .SP(n31694), .CK(debug_c_c), .Q(n1009));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D sub_62_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27242), 
          .S0(n931[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_9.INIT1 = 16'h0000;
    defparam sub_62_add_2_9.INJECT1_0 = "NO";
    defparam sub_62_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_62_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27241), 
          .COUT(n27242), .S0(n931[5]), .S1(n931[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_62_add_2_7.INJECT1_0 = "NO";
    defparam sub_62_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_62_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27240), 
          .COUT(n27241), .S0(n931[3]), .S1(n931[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_62_add_2_5.INJECT1_0 = "NO";
    defparam sub_62_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_62_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27239), 
          .COUT(n27240), .S0(n931[1]), .S1(n931[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_62_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_62_add_2_3.INJECT1_0 = "NO";
    defparam sub_62_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_62_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27239), 
          .S1(n931[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_62_add_2_1.INIT0 = 16'hF000;
    defparam sub_62_add_2_1.INIT1 = 16'h5555;
    defparam sub_62_add_2_1.INJECT1_0 = "NO";
    defparam sub_62_add_2_1.INJECT1_1 = "NO";
    LUT4 i15689_3_lut_rep_449 (.A(n27970), .B(n31789), .C(count[9]), .Z(n33442)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15689_3_lut_rep_449.init = 16'hecec;
    LUT4 i23213_3_lut_4_lut_4_lut (.A(n31740), .B(n33442), .C(n31731), 
         .D(n29512), .Z(n29778)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i23213_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i1_4_lut_adj_246 (.A(count[4]), .B(n29511), .C(count[3]), .D(n6), 
         .Z(n29512)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_246.init = 16'hccc8;
    LUT4 i21_3_lut_rep_307_4_lut_4_lut (.A(n27970), .B(n31789), .C(count[9]), 
         .D(n28201), .Z(n31730)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i21_3_lut_rep_307_4_lut_4_lut.init = 16'h1310;
    LUT4 i1_4_lut_adj_247 (.A(n31766), .B(count[8]), .C(n31851), .D(n31811), 
         .Z(n29416)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_247.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(count[4]), .B(n29381), .C(count[8]), .D(n29511), 
         .Z(n28201)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i22717_2_lut (.A(n1009), .B(n1021), .Z(n29864)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22717_2_lut.init = 16'hdddd;
    LUT4 i3_4_lut_adj_248 (.A(n28061), .B(n6_adj_183), .C(count[8]), .D(n31852), 
         .Z(n27970)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_248.init = 16'hfefc;
    LUT4 i3_4_lut_adj_249 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n28061)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_249.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6_adj_183)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3AX valid_48 (.D(n29778), .SP(n27924), .CK(debug_c_c), .Q(n1015));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(n1009), .B(n1021), .Z(n5_adj_182)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n29759), .D(n4), 
         .Z(n28181)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_250 (.A(n31868), .B(count[9]), .C(n28007), .D(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_250.init = 16'heccc;
    LUT4 i2_4_lut_adj_251 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28007)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_251.init = 16'hfeee;
    LUT4 i3073_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3073_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n29759)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_252 (.A(count[7]), .B(count[6]), .C(n31852), 
         .D(n29381), .Z(n29697)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_252.init = 16'h8000;
    LUT4 i3_3_lut_rep_366_4_lut (.A(count[12]), .B(n31869), .C(n29759), 
         .D(count[13]), .Z(n31789)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_366_4_lut.init = 16'hfffe;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    CCU2D add_1728_17 (.A0(count[15]), .B0(n5_adj_182), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26982), .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_17.INIT0 = 16'hd222;
    defparam add_1728_17.INIT1 = 16'h0000;
    defparam add_1728_17.INJECT1_0 = "NO";
    defparam add_1728_17.INJECT1_1 = "NO";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1728_15 (.A0(count[13]), .B0(n5_adj_182), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n5_adj_182), .C1(GND_net), 
          .D1(GND_net), .CIN(n26981), .COUT(n26982), .S0(n116[13]), 
          .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_15.INIT0 = 16'hd222;
    defparam add_1728_15.INIT1 = 16'hd222;
    defparam add_1728_15.INJECT1_0 = "NO";
    defparam add_1728_15.INJECT1_1 = "NO";
    CCU2D add_1728_13 (.A0(count[11]), .B0(n5_adj_182), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n5_adj_182), .C1(GND_net), 
          .D1(GND_net), .CIN(n26980), .COUT(n26981), .S0(n116[11]), 
          .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_13.INIT0 = 16'hd222;
    defparam add_1728_13.INIT1 = 16'hd222;
    defparam add_1728_13.INJECT1_0 = "NO";
    defparam add_1728_13.INJECT1_1 = "NO";
    CCU2D add_1728_11 (.A0(count[9]), .B0(n5_adj_182), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5_adj_182), .C1(GND_net), .D1(GND_net), 
          .CIN(n26979), .COUT(n26980), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_11.INIT0 = 16'hd222;
    defparam add_1728_11.INIT1 = 16'hd222;
    defparam add_1728_11.INJECT1_0 = "NO";
    defparam add_1728_11.INJECT1_1 = "NO";
    CCU2D add_1728_9 (.A0(count[7]), .B0(n5_adj_182), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5_adj_182), .C1(GND_net), .D1(GND_net), 
          .CIN(n26978), .COUT(n26979), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_9.INIT0 = 16'hd222;
    defparam add_1728_9.INIT1 = 16'hd222;
    defparam add_1728_9.INJECT1_0 = "NO";
    defparam add_1728_9.INJECT1_1 = "NO";
    CCU2D add_1728_7 (.A0(count[5]), .B0(n5_adj_182), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5_adj_182), .C1(GND_net), .D1(GND_net), 
          .CIN(n26977), .COUT(n26978), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_7.INIT0 = 16'hd222;
    defparam add_1728_7.INIT1 = 16'hd222;
    defparam add_1728_7.INJECT1_0 = "NO";
    defparam add_1728_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_253 (.A(n29416), .B(n931[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_253.init = 16'h4444;
    CCU2D add_1728_5 (.A0(count[3]), .B0(n5_adj_182), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5_adj_182), .C1(GND_net), .D1(GND_net), 
          .CIN(n26976), .COUT(n26977), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1728_5.INIT0 = 16'hd222;
    defparam add_1728_5.INIT1 = 16'hd222;
    defparam add_1728_5.INJECT1_0 = "NO";
    defparam add_1728_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_308_3_lut (.A(count[9]), .B(n31789), .C(count[8]), 
         .Z(n31731)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_308_3_lut.init = 16'hfefe;
    LUT4 i23134_4_lut (.A(n31730), .B(n29864), .C(n29416), .D(n10), 
         .Z(n30189)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23134_4_lut.init = 16'h3323;
    LUT4 i8_4_lut (.A(n31812), .B(n16), .C(count[13]), .D(count[11]), 
         .Z(n16124)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i8_4_lut.init = 16'h0004;
    LUT4 i7_4_lut (.A(count[10]), .B(n31694), .C(n26), .D(n29864), .Z(n16)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i7_4_lut.init = 16'h0040;
    LUT4 i33_3_lut (.A(n28201), .B(n27970), .C(count[9]), .Z(n26)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut_adj_254 (.A(n29416), .B(n931[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_254.init = 16'h4444;
    LUT4 i1_2_lut_adj_255 (.A(n29416), .B(n931[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_255.init = 16'h4444;
    LUT4 i1_2_lut_adj_256 (.A(n29416), .B(n931[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_256.init = 16'h4444;
    LUT4 i1_2_lut_adj_257 (.A(n29416), .B(n931[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_257.init = 16'h4444;
    LUT4 i1_2_lut_adj_258 (.A(n29416), .B(n931[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_258.init = 16'h4444;
    LUT4 i1_2_lut_adj_259 (.A(n29416), .B(n931[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_259.init = 16'h4444;
    LUT4 i1_2_lut_adj_260 (.A(n29416), .B(n931[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_260.init = 16'h4444;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14183), .PD(n16124), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (n30186, GND_net, debug_c_c, n31694, rc_ch2_c, 
            n1000, n27915, \register[2] , n14186, n30218) /* synthesis syn_module_defined=1 */ ;
    output n30186;
    input GND_net;
    input debug_c_c;
    input n31694;
    input rc_ch2_c;
    output n1000;
    input n27915;
    output [7:0]\register[2] ;
    input n14186;
    output n30218;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n1006, n994, n31862, n28054, n31863, n31738, n29784;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31864, n28047, n5, n31865, n28046, n27833, n31866, n29688, 
        n29920, n31792, n31769, n27246;
    wire [7:0]n922;
    
    wire n27245, n27244, n31793, n22003, n13322, n27243, n31770, 
        n31771, n31737, n29785, n29934, n29974, n13384, n29770, 
        n26990;
    wire [15:0]n116;
    
    wire n26989, n26988, n26987, n26986, n26985, n26984, n26983, 
        n16127;
    wire [7:0]n43;
    
    wire n29678, n29768, n4, n6, n29469, n31736;
    
    LUT4 i1_2_lut_rep_439 (.A(n1006), .B(n994), .Z(n31862)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_439.init = 16'hbbbb;
    LUT4 i23131_2_lut_3_lut (.A(n1006), .B(n994), .C(n28054), .Z(n30186)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i23131_2_lut_3_lut.init = 16'h4040;
    LUT4 i5_2_lut_rep_440 (.A(n994), .B(n1006), .Z(n31863)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_440.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n994), .B(n1006), .C(n31738), .Z(n29784)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_rep_441 (.A(count[4]), .B(count[5]), .Z(n31864)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_441.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(n28047), .D(count[6]), 
         .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_442 (.A(count[7]), .B(count[6]), .Z(n31865)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_442.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n28046), .D(count[5]), 
         .Z(n27833)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_443 (.A(count[2]), .B(count[3]), .Z(n31866)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_443.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_237 (.A(count[2]), .B(count[3]), .C(count[1]), 
         .Z(n29688)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_adj_237.init = 16'h8080;
    LUT4 i2_2_lut_rep_369 (.A(count[0]), .B(n29920), .Z(n31792)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_rep_369.init = 16'h8888;
    LUT4 i1_2_lut_rep_346_3_lut (.A(count[0]), .B(n29920), .C(count[8]), 
         .Z(n31769)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_346_3_lut.init = 16'h8080;
    CCU2D sub_61_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27246), 
          .S0(n922[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_61_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_9.INIT1 = 16'h0000;
    defparam sub_61_add_2_9.INJECT1_0 = "NO";
    defparam sub_61_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27245), 
          .COUT(n27246), .S0(n922[5]), .S1(n922[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_61_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_7.INJECT1_0 = "NO";
    defparam sub_61_add_2_7.INJECT1_1 = "NO";
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n31694), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1006));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    CCU2D sub_61_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27244), 
          .COUT(n27245), .S0(n922[3]), .S1(n922[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_61_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_5.INJECT1_0 = "NO";
    defparam sub_61_add_2_5.INJECT1_1 = "NO";
    LUT4 i15620_2_lut_3_lut_4_lut (.A(count[0]), .B(n29920), .C(n31793), 
         .D(count[8]), .Z(n22003)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i15620_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_370 (.A(count[9]), .B(n13322), .Z(n31793)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_370.init = 16'heeee;
    CCU2D sub_61_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27243), 
          .COUT(n27244), .S0(n922[1]), .S1(n922[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_61_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_3.INJECT1_0 = "NO";
    defparam sub_61_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27243), 
          .S1(n922[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_61_add_2_1.INIT0 = 16'hF000;
    defparam sub_61_add_2_1.INIT1 = 16'h5555;
    defparam sub_61_add_2_1.INJECT1_0 = "NO";
    defparam sub_61_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_347_4_lut (.A(count[9]), .B(n13322), .C(n29920), 
         .D(count[8]), .Z(n31770)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_3_lut_rep_347_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_348_3_lut (.A(count[9]), .B(n13322), .C(count[8]), 
         .Z(n31771)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_348_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_314_3_lut_4_lut (.A(count[9]), .B(n13322), .C(n27833), 
         .D(count[8]), .Z(n31737)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_314_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX valid_48 (.D(n29785), .SP(n27915), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1000));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i22822_3_lut_4_lut (.A(n31769), .B(n29934), .C(n31793), .D(n31770), 
         .Z(n29974)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i22822_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23186_3_lut_3_lut_4_lut (.A(n27833), .B(n31771), .C(n29934), 
         .D(n31738), .Z(n29785)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23186_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i22673_4_lut_rep_315 (.A(n13384), .B(count[13]), .C(count[12]), 
         .D(n29770), .Z(n31738)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i22673_4_lut_rep_315.init = 16'heaaa;
    CCU2D add_1724_17 (.A0(count[15]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26990), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_17.INIT0 = 16'hd222;
    defparam add_1724_17.INIT1 = 16'h0000;
    defparam add_1724_17.INJECT1_0 = "NO";
    defparam add_1724_17.INJECT1_1 = "NO";
    CCU2D add_1724_15 (.A0(count[13]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31863), .C1(GND_net), .D1(GND_net), .CIN(n26989), 
          .COUT(n26990), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_15.INIT0 = 16'hd222;
    defparam add_1724_15.INIT1 = 16'hd222;
    defparam add_1724_15.INJECT1_0 = "NO";
    defparam add_1724_15.INJECT1_1 = "NO";
    CCU2D add_1724_13 (.A0(count[11]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31863), .C1(GND_net), .D1(GND_net), .CIN(n26988), 
          .COUT(n26989), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_13.INIT0 = 16'hd222;
    defparam add_1724_13.INIT1 = 16'hd222;
    defparam add_1724_13.INJECT1_0 = "NO";
    defparam add_1724_13.INJECT1_1 = "NO";
    CCU2D add_1724_11 (.A0(count[9]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31863), .C1(GND_net), .D1(GND_net), .CIN(n26987), 
          .COUT(n26988), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_11.INIT0 = 16'hd222;
    defparam add_1724_11.INIT1 = 16'hd222;
    defparam add_1724_11.INJECT1_0 = "NO";
    defparam add_1724_11.INJECT1_1 = "NO";
    CCU2D add_1724_9 (.A0(count[7]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31863), .C1(GND_net), .D1(GND_net), .CIN(n26986), 
          .COUT(n26987), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_9.INIT0 = 16'hd222;
    defparam add_1724_9.INIT1 = 16'hd222;
    defparam add_1724_9.INJECT1_0 = "NO";
    defparam add_1724_9.INJECT1_1 = "NO";
    CCU2D add_1724_7 (.A0(count[5]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31863), .C1(GND_net), .D1(GND_net), .CIN(n26985), 
          .COUT(n26986), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_7.INIT0 = 16'hd222;
    defparam add_1724_7.INIT1 = 16'hd222;
    defparam add_1724_7.INJECT1_0 = "NO";
    defparam add_1724_7.INJECT1_1 = "NO";
    CCU2D add_1724_5 (.A0(count[3]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31863), .C1(GND_net), .D1(GND_net), .CIN(n26984), 
          .COUT(n26985), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_5.INIT0 = 16'hd222;
    defparam add_1724_5.INIT1 = 16'hd222;
    defparam add_1724_5.INJECT1_0 = "NO";
    defparam add_1724_5.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    CCU2D add_1724_3 (.A0(count[1]), .B0(n31863), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31863), .C1(GND_net), .D1(GND_net), .CIN(n26983), 
          .COUT(n26984), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_3.INIT0 = 16'hd222;
    defparam add_1724_3.INIT1 = 16'hd222;
    defparam add_1724_3.INJECT1_0 = "NO";
    defparam add_1724_3.INJECT1_1 = "NO";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    CCU2D add_1724_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29784), .B1(n1006), .C1(count[0]), .D1(n994), .COUT(n26983), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1724_1.INIT0 = 16'hF000;
    defparam add_1724_1.INIT1 = 16'ha565;
    defparam add_1724_1.INJECT1_0 = "NO";
    defparam add_1724_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1006), .SP(n31694), .CK(debug_c_c), .Q(n994));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i23163_4_lut (.A(n29678), .B(n31863), .C(n31738), .D(n31862), 
         .Z(n30218)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i23163_4_lut.init = 16'h3031;
    LUT4 i3_4_lut (.A(n31771), .B(n29974), .C(n31792), .D(n27833), .Z(n29678)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut.init = 16'h3222;
    LUT4 i2_4_lut (.A(n29768), .B(count[9]), .C(count[8]), .D(n4), .Z(n29770)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut.init = 16'hfeee;
    LUT4 i1_4_lut (.A(n31865), .B(count[4]), .C(count[5]), .D(n29688), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut.init = 16'haaa8;
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n29768)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i22785_4_lut (.A(n13322), .B(count[9]), .C(n5), .D(n6), .Z(n29934)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i22785_4_lut.init = 16'heeea;
    LUT4 i2_2_lut (.A(count[7]), .B(count[8]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_238 (.A(count[2]), .B(count[1]), .C(count[0]), .D(count[3]), 
         .Z(n28047)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_4_lut_adj_238.init = 16'hfffe;
    LUT4 i3_4_lut_adj_239 (.A(count[12]), .B(count[13]), .C(n13384), .D(n29768), 
         .Z(n13322)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_239.init = 16'hfffe;
    LUT4 i1_2_lut_adj_240 (.A(count[15]), .B(count[14]), .Z(n13384)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_240.init = 16'heeee;
    LUT4 i2_4_lut_adj_241 (.A(count[2]), .B(count[4]), .C(count[1]), .D(count[3]), 
         .Z(n28046)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_241.init = 16'hffec;
    LUT4 i22773_4_lut (.A(count[1]), .B(n31866), .C(n31865), .D(n31864), 
         .Z(n29920)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22773_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_242 (.A(n994), .B(n31694), .C(n29469), .D(n29934), 
         .Z(n16127)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_242.init = 16'h0080;
    LUT4 i2_4_lut_adj_243 (.A(n31769), .B(n28054), .C(count[9]), .D(n1006), 
         .Z(n29469)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_243.init = 16'h00c8;
    LUT4 i2_4_lut_adj_244 (.A(n31736), .B(n31770), .C(n31737), .D(n22003), 
         .Z(n28054)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_244.init = 16'heefe;
    LUT4 i21_3_lut_rep_313_4_lut (.A(count[8]), .B(n31792), .C(n31793), 
         .D(n29934), .Z(n31736)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21_3_lut_rep_313_4_lut.init = 16'h00f8;
    LUT4 i15334_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15334_2_lut_4_lut.init = 16'h0200;
    LUT4 i15333_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15333_2_lut_4_lut.init = 16'h0200;
    LUT4 i15332_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15332_2_lut_4_lut.init = 16'h0200;
    LUT4 i15331_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15331_2_lut_4_lut.init = 16'h0200;
    LUT4 i15330_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15330_2_lut_4_lut.init = 16'h0200;
    LUT4 i15329_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15329_2_lut_4_lut.init = 16'h0200;
    LUT4 i15328_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15328_2_lut_4_lut.init = 16'h0200;
    LUT4 i15089_2_lut_4_lut (.A(count[8]), .B(n31793), .C(n29920), .D(n922[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15089_2_lut_4_lut.init = 16'h0200;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14186), .PD(n16127), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (GND_net, debug_c_c, n31694, n29930, \register[1] , 
            n14187, n9, rc_ch1_c, n30152, n30184, n985, n27912) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n31694;
    output n29930;
    output [7:0]\register[1] ;
    input n14187;
    input n9;
    input rc_ch1_c;
    output n30152;
    output n30184;
    output n985;
    input n27912;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n979, n991, n31853, n31756, n29787;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n13308, n31782, n31753, n31755, n21922, n29637, n31725, 
        n27250;
    wire [7:0]n913;
    
    wire n27249, n27248, n27247, n31726, n23, n29976;
    wire [15:0]n116;
    
    wire n26998, n26997, n26996, n26995, n26994, n26993, n26992, 
        n26991, n16131;
    wire [7:0]n43;
    
    wire n29762, n28038, n4, n29764, n6, n13393, n28093, n8, 
        n95, n49_adj_181, n30027, n29978, n29635, n31714, n29681, 
        n31839, n29788;
    
    LUT4 i5_2_lut_rep_430 (.A(n979), .B(n991), .Z(n31853)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_430.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n979), .B(n991), .C(n31756), .Z(n29787)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_rep_359 (.A(count[9]), .B(n13308), .Z(n31782)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_359.init = 16'heeee;
    LUT4 i1_2_lut_rep_330_3_lut (.A(count[9]), .B(n13308), .C(count[8]), 
         .Z(n31753)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_330_3_lut.init = 16'hfefe;
    LUT4 i15542_2_lut_3_lut_4_lut (.A(count[9]), .B(n13308), .C(n31755), 
         .D(count[8]), .Z(n21922)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i15542_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_302_3_lut_4_lut (.A(count[9]), .B(n13308), .C(n29637), 
         .D(count[8]), .Z(n31725)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_302_3_lut_4_lut.init = 16'hfffe;
    CCU2D sub_60_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27250), 
          .S0(n913[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_60_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_9.INIT1 = 16'h0000;
    defparam sub_60_add_2_9.INJECT1_0 = "NO";
    defparam sub_60_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27249), 
          .COUT(n27250), .S0(n913[5]), .S1(n913[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_60_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_7.INJECT1_0 = "NO";
    defparam sub_60_add_2_7.INJECT1_1 = "NO";
    FD1P3AX prev_in_46 (.D(n991), .SP(n31694), .CK(debug_c_c), .Q(n979));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D sub_60_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27248), 
          .COUT(n27249), .S0(n913[3]), .S1(n913[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_60_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_5.INJECT1_0 = "NO";
    defparam sub_60_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27247), 
          .COUT(n27248), .S0(n913[1]), .S1(n913[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_60_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_3.INJECT1_0 = "NO";
    defparam sub_60_add_2_3.INJECT1_1 = "NO";
    LUT4 i22824_3_lut_4_lut (.A(n31726), .B(n29930), .C(n31782), .D(n23), 
         .Z(n29976)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i22824_3_lut_4_lut.init = 16'hfffe;
    CCU2D sub_60_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27247), 
          .S1(n913[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_60_add_2_1.INIT0 = 16'hF000;
    defparam sub_60_add_2_1.INIT1 = 16'h5555;
    defparam sub_60_add_2_1.INJECT1_0 = "NO";
    defparam sub_60_add_2_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    CCU2D add_1720_17 (.A0(count[15]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26998), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_17.INIT0 = 16'hd222;
    defparam add_1720_17.INIT1 = 16'h0000;
    defparam add_1720_17.INJECT1_0 = "NO";
    defparam add_1720_17.INJECT1_1 = "NO";
    CCU2D add_1720_15 (.A0(count[13]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31853), .C1(GND_net), .D1(GND_net), .CIN(n26997), 
          .COUT(n26998), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_15.INIT0 = 16'hd222;
    defparam add_1720_15.INIT1 = 16'hd222;
    defparam add_1720_15.INJECT1_0 = "NO";
    defparam add_1720_15.INJECT1_1 = "NO";
    CCU2D add_1720_13 (.A0(count[11]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31853), .C1(GND_net), .D1(GND_net), .CIN(n26996), 
          .COUT(n26997), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_13.INIT0 = 16'hd222;
    defparam add_1720_13.INIT1 = 16'hd222;
    defparam add_1720_13.INJECT1_0 = "NO";
    defparam add_1720_13.INJECT1_1 = "NO";
    CCU2D add_1720_11 (.A0(count[9]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31853), .C1(GND_net), .D1(GND_net), .CIN(n26995), 
          .COUT(n26996), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_11.INIT0 = 16'hd222;
    defparam add_1720_11.INIT1 = 16'hd222;
    defparam add_1720_11.INJECT1_0 = "NO";
    defparam add_1720_11.INJECT1_1 = "NO";
    CCU2D add_1720_9 (.A0(count[7]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31853), .C1(GND_net), .D1(GND_net), .CIN(n26994), 
          .COUT(n26995), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_9.INIT0 = 16'hd222;
    defparam add_1720_9.INIT1 = 16'hd222;
    defparam add_1720_9.INJECT1_0 = "NO";
    defparam add_1720_9.INJECT1_1 = "NO";
    CCU2D add_1720_7 (.A0(count[5]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31853), .C1(GND_net), .D1(GND_net), .CIN(n26993), 
          .COUT(n26994), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_7.INIT0 = 16'hd222;
    defparam add_1720_7.INIT1 = 16'hd222;
    defparam add_1720_7.INJECT1_0 = "NO";
    defparam add_1720_7.INJECT1_1 = "NO";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    CCU2D add_1720_5 (.A0(count[3]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31853), .C1(GND_net), .D1(GND_net), .CIN(n26992), 
          .COUT(n26993), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_5.INIT0 = 16'hd222;
    defparam add_1720_5.INIT1 = 16'hd222;
    defparam add_1720_5.INJECT1_0 = "NO";
    defparam add_1720_5.INJECT1_1 = "NO";
    CCU2D add_1720_3 (.A0(count[1]), .B0(n31853), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31853), .C1(GND_net), .D1(GND_net), .CIN(n26991), 
          .COUT(n26992), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_3.INIT0 = 16'hd222;
    defparam add_1720_3.INIT1 = 16'hd222;
    defparam add_1720_3.INJECT1_0 = "NO";
    defparam add_1720_3.INJECT1_1 = "NO";
    CCU2D add_1720_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29787), .B1(n991), .C1(count[0]), .D1(n979), .COUT(n26991), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1720_1.INIT0 = 16'hF000;
    defparam add_1720_1.INIT1 = 16'ha565;
    defparam add_1720_1.INJECT1_0 = "NO";
    defparam add_1720_1.INJECT1_1 = "NO";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n29762), .B(count[9]), .C(n28038), .D(n4), .Z(n29764)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut.init = 16'hfeee;
    LUT4 i2_4_lut_adj_229 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28038)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_229.init = 16'hfeee;
    LUT4 i3189_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3189_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n29762)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_230 (.A(count[15]), .B(count[14]), .Z(n13393)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_230.init = 16'heeee;
    LUT4 i5_4_lut (.A(n9), .B(n28093), .C(n8), .D(n979), .Z(n16131)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i15327_2_lut (.A(n913[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15327_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(count[8]), .B(n31782), .C(count[1]), .D(n95), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0222;
    LUT4 i22782_4_lut (.A(n13308), .B(count[9]), .C(n49_adj_181), .D(n30027), 
         .Z(n29930)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i22782_4_lut.init = 16'heeea;
    LUT4 i2_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n49_adj_181)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n31694), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n991));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i22874_4_lut (.A(count[4]), .B(count[1]), .C(count[5]), .D(n29978), 
         .Z(n30027)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i22874_4_lut.init = 16'ha080;
    LUT4 i22826_3_lut (.A(count[0]), .B(count[2]), .C(count[3]), .Z(n29978)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22826_3_lut.init = 16'hfefe;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n13393), .D(n29762), 
         .Z(n13308)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_231 (.A(count[3]), .B(count[4]), .C(count[2]), .D(n29635), 
         .Z(n95)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_231.init = 16'h8000;
    LUT4 i2_4_lut_adj_232 (.A(n31714), .B(n23), .C(n31725), .D(n21922), 
         .Z(n28093)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_232.init = 16'heefe;
    LUT4 i1_4_lut_adj_233 (.A(count[4]), .B(n29635), .C(count[3]), .D(n6), 
         .Z(n29637)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_233.init = 16'hccc8;
    LUT4 i15326_2_lut (.A(n913[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15326_2_lut.init = 16'h8888;
    LUT4 i23097_4_lut (.A(n29681), .B(n31853), .C(n31756), .D(n31839), 
         .Z(n30152)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i23097_4_lut.init = 16'h3031;
    LUT4 i3_4_lut_adj_234 (.A(n31753), .B(n29976), .C(n31755), .D(n29637), 
         .Z(n29681)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut_adj_234.init = 16'h3222;
    LUT4 i15325_2_lut (.A(n913[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15325_2_lut.init = 16'h8888;
    LUT4 i15324_2_lut (.A(n913[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15324_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_416 (.A(n991), .B(n979), .Z(n31839)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_416.init = 16'hbbbb;
    LUT4 i23129_2_lut_3_lut (.A(n991), .B(n979), .C(n28093), .Z(n30184)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i23129_2_lut_3_lut.init = 16'h4040;
    LUT4 i23184_3_lut_3_lut_4_lut (.A(n29637), .B(n31753), .C(n29930), 
         .D(n31756), .Z(n29788)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23184_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i21_3_lut_rep_291_4_lut (.A(count[8]), .B(n31755), .C(n31782), 
         .D(n29930), .Z(n31714)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21_3_lut_rep_291_4_lut.init = 16'h00f8;
    LUT4 i2_3_lut_4_lut (.A(count[8]), .B(n31755), .C(count[9]), .D(n991), 
         .Z(n8)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_3_lut_4_lut.init = 16'h00f8;
    LUT4 i1_2_lut_3_lut_adj_235 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_adj_235.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_236 (.A(count[6]), .B(count[7]), .C(count[5]), 
         .Z(n29635)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_adj_236.init = 16'h8080;
    LUT4 i15084_2_lut (.A(n913[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15084_2_lut.init = 16'h8888;
    LUT4 i15323_2_lut (.A(n913[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15323_2_lut.init = 16'h8888;
    LUT4 i15322_2_lut (.A(n913[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15322_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_rep_332 (.A(n95), .B(count[1]), .C(count[0]), .Z(n31755)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_332.init = 16'h8080;
    LUT4 i1_2_lut_rep_303_4_lut (.A(n95), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n31726)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_303_4_lut.init = 16'h8000;
    LUT4 i15321_2_lut (.A(n913[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15321_2_lut.init = 16'h8888;
    LUT4 i22761_4_lut_rep_333 (.A(n13393), .B(count[13]), .C(count[12]), 
         .D(n29764), .Z(n31756)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i22761_4_lut_rep_333.init = 16'heaaa;
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX valid_48 (.D(n29788), .SP(n27912), .CD(GND_net), .CK(debug_c_c), 
            .Q(n985));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14187), .PD(n16131), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n31694), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n31694), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (debug_c_c, n33455, \select[7] , 
            \select[1] , \select[4] , \select[2] , databus_out, n13568, 
            \read_value[6] , n33446, n2, register_addr, n31751, \read_value[3] , 
            rw, n2_adj_43, \register[2][0] , \register_addr[3] , n31716, 
            \register_addr[1] , \steps_reg[5] , n14, \read_value[4] , 
            n2_adj_44, n31827, n27707, n31720, n33447, n14124, \read_value[7] , 
            n2_adj_45, n1306, \read_value[2] , n2_adj_46, n1309, n1312, 
            \read_value[1] , n2_adj_47, \read_value[0] , n2_adj_48, 
            \read_value[5] , n2_adj_49, n31717, n31867, n31698, n191, 
            n29590, n31699, n13671, n31705, n8940, \sendcount[1] , 
            prev_select, n2658, n21, n29452, n185, n14252, \register_addr[4] , 
            n31746, debug_c_7, n13757, n31779, n29552, n47, \read_size[2] , 
            n6, n31739, \read_value[1]_adj_50 , n4, n3970, n78, 
            n31763, \read_value[19] , n3, \read_value[20] , n3_adj_51, 
            \read_size[2]_adj_52 , n31832, \read_value[21] , n3_adj_53, 
            prev_select_adj_54, n14172, \read_value[22] , n3_adj_55, 
            \read_value[23] , n3_adj_56, \read_value[24] , n3_adj_57, 
            \read_value[25] , n3_adj_58, \read_value[26] , n3_adj_59, 
            \read_value[27] , n3_adj_60, \read_value[28] , n3_adj_61, 
            \read_value[29] , n3_adj_62, \read_value[30] , n3_adj_63, 
            n31741, \read_value[31] , n3_adj_64, \read_value[18] , n3_adj_65, 
            \read_value[17] , n3_adj_66, \read_value[16] , n3_adj_67, 
            \read_value[15] , n3_adj_68, \read_value[14] , n3_adj_69, 
            \read_value[13] , n3_adj_70, n31783, databus, \read_value[12] , 
            n3_adj_71, \read_value[11] , n3_adj_72, \read_value[10] , 
            n3_adj_73, n28025, n33445, n33457, n28937, n31780, \read_value[9] , 
            n3_adj_74, n22093, \read_value[8] , n3_adj_75, n31762, 
            prev_select_adj_76, n29823, n31703, n31718, n31774, n14022, 
            n16046, n16045, n24748, n250, \read_value[1]_adj_77 , 
            n1, n29738, \steps_reg[6] , n13, n31724, n12795, n9, 
            n14_adj_78, n10, \reg_size[2] , n31841, n106, \control_reg[7] , 
            n8243, \read_size[0] , \read_size[0]_adj_79 , n55, \read_size[2]_adj_80 , 
            n9_adj_81, \control_reg[7]_adj_82 , n1_adj_83, n5613, n31722, 
            n13779, n31707, n31785, n14084, \read_size[0]_adj_84 , 
            n29694, n13476, \control_reg[7]_adj_85 , n8252, n4_adj_86, 
            \control_reg[7]_adj_87 , n8261, n31733, \steps_reg[3] , 
            n12, \arm_select[0] , n31727, prev_select_adj_88, n3883, 
            n9089, n24720, n24690, n13606, n89, n31732, n3786, 
            n31700, n3700, n8885, debug_c_2, debug_c_3, debug_c_4, 
            debug_c_5, n31701, n24729, n31708, prev_select_adj_89, 
            n31715, n31719, n10607, GND_net, n10608_c) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n33455;
    output \select[7] ;
    output \select[1] ;
    output \select[4] ;
    output \select[2] ;
    output [31:0]databus_out;
    input n13568;
    input \read_value[6] ;
    output n33446;
    output n2;
    output [7:0]register_addr;
    input n31751;
    input \read_value[3] ;
    output rw;
    output n2_adj_43;
    input \register[2][0] ;
    output \register_addr[3] ;
    output n31716;
    output \register_addr[1] ;
    input \steps_reg[5] ;
    output n14;
    input \read_value[4] ;
    output n2_adj_44;
    output n31827;
    output n27707;
    output n31720;
    input n33447;
    output n14124;
    input \read_value[7] ;
    output n2_adj_45;
    output n1306;
    input \read_value[2] ;
    output n2_adj_46;
    output n1309;
    output n1312;
    input \read_value[1] ;
    output n2_adj_47;
    input \read_value[0] ;
    output n2_adj_48;
    input \read_value[5] ;
    output n2_adj_49;
    output n31717;
    input n31867;
    output n31698;
    output n191;
    output n29590;
    output n31699;
    input n13671;
    output n31705;
    output n8940;
    output \sendcount[1] ;
    input prev_select;
    output n2658;
    input n21;
    output n29452;
    input n185;
    output n14252;
    output \register_addr[4] ;
    output n31746;
    output debug_c_7;
    output n13757;
    output n31779;
    output n29552;
    output n47;
    input \read_size[2] ;
    output n6;
    output n31739;
    input \read_value[1]_adj_50 ;
    output n4;
    output n3970;
    output n78;
    output n31763;
    input \read_value[19] ;
    output n3;
    input \read_value[20] ;
    output n3_adj_51;
    input \read_size[2]_adj_52 ;
    input n31832;
    input \read_value[21] ;
    output n3_adj_53;
    input prev_select_adj_54;
    output n14172;
    input \read_value[22] ;
    output n3_adj_55;
    input \read_value[23] ;
    output n3_adj_56;
    input \read_value[24] ;
    output n3_adj_57;
    input \read_value[25] ;
    output n3_adj_58;
    input \read_value[26] ;
    output n3_adj_59;
    input \read_value[27] ;
    output n3_adj_60;
    input \read_value[28] ;
    output n3_adj_61;
    input \read_value[29] ;
    output n3_adj_62;
    input \read_value[30] ;
    output n3_adj_63;
    output n31741;
    input \read_value[31] ;
    output n3_adj_64;
    input \read_value[18] ;
    output n3_adj_65;
    input \read_value[17] ;
    output n3_adj_66;
    input \read_value[16] ;
    output n3_adj_67;
    input \read_value[15] ;
    output n3_adj_68;
    input \read_value[14] ;
    output n3_adj_69;
    input \read_value[13] ;
    output n3_adj_70;
    input n31783;
    input [31:0]databus;
    input \read_value[12] ;
    output n3_adj_71;
    input \read_value[11] ;
    output n3_adj_72;
    input \read_value[10] ;
    output n3_adj_73;
    input n28025;
    input n33445;
    output n33457;
    output n28937;
    output n31780;
    input \read_value[9] ;
    output n3_adj_74;
    output n22093;
    input \read_value[8] ;
    output n3_adj_75;
    output n31762;
    input prev_select_adj_76;
    output n29823;
    output n31703;
    output n31718;
    output n31774;
    input n14022;
    output n16046;
    output n16045;
    output n24748;
    output n250;
    input \read_value[1]_adj_77 ;
    output n1;
    output n29738;
    input \steps_reg[6] ;
    output n13;
    output n31724;
    input n12795;
    input n9;
    input n14_adj_78;
    input n10;
    input \reg_size[2] ;
    input n31841;
    output n106;
    input \control_reg[7] ;
    output n8243;
    input \read_size[0] ;
    input \read_size[0]_adj_79 ;
    output n55;
    input \read_size[2]_adj_80 ;
    output n9_adj_81;
    input \control_reg[7]_adj_82 ;
    output n1_adj_83;
    output n5613;
    output n31722;
    output n13779;
    output n31707;
    output n31785;
    output n14084;
    input \read_size[0]_adj_84 ;
    output n29694;
    output n13476;
    input \control_reg[7]_adj_85 ;
    output n8252;
    output n4_adj_86;
    input \control_reg[7]_adj_87 ;
    output n8261;
    output n31733;
    input \steps_reg[3] ;
    output n12;
    output \arm_select[0] ;
    output n31727;
    input prev_select_adj_88;
    output n3883;
    output n9089;
    output n24720;
    output n24690;
    output n13606;
    output n89;
    output n31732;
    output n3786;
    output n31700;
    output n3700;
    output n8885;
    output debug_c_2;
    output debug_c_3;
    output debug_c_4;
    output debug_c_5;
    output n31701;
    output n24729;
    output n31708;
    input prev_select_adj_89;
    output n31715;
    output n31719;
    output n10607;
    input GND_net;
    input n10608_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire n33445 /* synthesis nomerge= */ ;
    wire n31780 /* synthesis SET_AS_NETWORK=n31780 */ ;
    wire n31762 /* synthesis SET_AS_NETWORK=n31762 */ ;
    wire [31:0]n1294;
    
    wire n1747;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n31757;
    wire [4:0]n18;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n12_c, n13456, n15880, n15875, n29263;
    wire [127:0]select;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    
    wire n31686, n15886, n31687, n2619;
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n29640;
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n15879;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n31750;
    wire [7:0]n2036;
    
    wire n15885;
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n15872;
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    
    wire n30802;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n30672, n29639;
    wire [7:0]n5604;
    
    wire n31765, n2617;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n31887, n33438, n15046, n21320, n28985, n29956, n29428;
    wire [7:0]register_addr_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire n11867, n10734, n29123, n11865, n10743, n1406, n1405, 
        n1399, n29655, n29418, n11698, n29153, n29187, n31728, 
        n31236, n29708, n29709;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n29632, n31807, n31822, n31874, n31873, n31877, n31876;
    wire [4:0]n19;
    
    wire n31745, n29623, n31806, n31880, n31879, n4_c, n31723, 
        n29710, n31883, escape, n31238, n31882, n31886, n31885, 
        n31889, n31888, n29419, n15, n30012, n13070, n29758, n31892, 
        n31795, n13182, n8, n31891, n31901, n31900, n31904, n31903, 
        n32225, n29699, n160, n10514, n29757, n31754, n20, n29808, 
        n9_adj_74, n31830, n2045, n31706, n11_adj_81, n14_adj_82, 
        n28977, n30796, n11_adj_83, n28981, n11_adj_85, n28983, 
        n11_adj_87, n28991, n32223, n11_adj_89, n28989, n11_adj_91, 
        n28987, n11_adj_92, n29059, n11_adj_96, n28979, n31815, 
        n11_adj_99, n11_adj_102, n28959, n6_adj_103, n11_adj_104, 
        n29039, n11_adj_106, n29055, n11_adj_107, n29095, n11_adj_108, 
        n29047, n11_adj_109, n29011, n11_adj_110, n28969, n5, n29523, 
        n28079, n31829, n31805, n4_adj_111, n31893;
    wire [7:0]n9241;
    
    wire n5_adj_112, n29532, n28074, n5_adj_113, n29522, n28077, 
        n4_adj_116, n31881, send, n4_adj_118, n31875, n31787, n31828, 
        n31817, n31781, n28097, n31834, n31890, n30800, n30801, 
        n31871, n4_adj_119, n31902, n4_adj_120, n31905, n4_adj_121, 
        n31872, n4_adj_122, n31878, n15_adj_123, n31840, n5_adj_124, 
        n29524, n28075, n5_adj_127, n29525, n28076, n5_adj_128, 
        n29526, n28072, n5_adj_130, n29527, n28091, n31772, n5_adj_131, 
        n29528, n28073, n5_adj_132, n29529, n28034, n30673, n29767, 
        n29766, n28151, n29744, n5_adj_133, n29531, n28086, n5_adj_134, 
        n29521, n27895, n5_adj_135, n29516, n28005, n5_adj_136, 
        n29534, n28083, n31870, n16067, n31816, n30016, n5_adj_137, 
        n29530, n28022, n31804, n31235, n7, n5_adj_139, n29519, 
        n28008, n5_adj_140, n29536, n28084, n5_adj_141, n29535, 
        n28082, n2557, n31823, n29795, n31824, n15045;
    wire [3:0]n1690;
    
    wire n1695, n31825, n9_adj_142, n8_adj_143, n15871, n6_adj_144, 
        n5_adj_145, n29533, n28048, n31826, n29874, n1_adj_147, 
        n6_adj_148, n29404, n5_adj_151, n29537, n28035, n5_adj_155, 
        n29538, n28002, n9017, n5_adj_158, n29539, n28016, n27964, 
        n28012, n28030, n27994, n27999, n28013, n28023, n28026, 
        n27998, n28020, n28019, n5_adj_159, n29540, n5_adj_160, 
        n29541, n5_adj_161, n29542, n31833, n30674, n5_adj_162, 
        n29543;
    wire [3:0]n17;
    
    wire n16049, n5_adj_163, n29544, n5_adj_164, n29545, n5_adj_165, 
        n29546, n5_adj_166, n29515, n5_adj_167, n29520, n31794, 
        n5_adj_168, n29517, busy, n29627, n5_adj_170, n29518, n29860, 
        n30831, n29912, n21052, n29980, n29473, n38, n31773, n4_adj_176, 
        n8_adj_177, n4_adj_178, n6_adj_179;
    
    LUT4 i1_2_lut (.A(n1294[6]), .B(n1294[11]), .Z(n1747)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3AX sendcount__i0 (.D(n18[0]), .SP(n31757), .CK(debug_c_c), .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(\buffer[0] [3]), .B(\buffer[0] [5]), .C(\buffer[0] [4]), 
         .D(\buffer[0] [6]), .Z(n12_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i3_4_lut.init = 16'hfffe;
    FD1S3JX state_FSM_i1 (.D(n13456), .CK(debug_c_c), .PD(n33455), .Q(n1294[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1S3IX select__i7 (.D(n15880), .CK(debug_c_c), .CD(n33455), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 i15447_2_lut_3_lut (.A(n1294[0]), .B(n1294[8]), .C(\select[1] ), 
         .Z(n15875)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15447_2_lut_3_lut.init = 16'h1010;
    FD1S3IX select__i4 (.D(n29263), .CK(debug_c_c), .CD(n33455), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1S3IX select__i3 (.D(n31686), .CK(debug_c_c), .CD(n33455), .Q(select[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i3.GSR = "ENABLED";
    FD1S3IX select__i2 (.D(n15886), .CK(debug_c_c), .CD(n33455), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1S3IX select__i1 (.D(n31687), .CK(debug_c_c), .CD(n33455), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(n1294[0]), .B(n1294[8]), .C(select[3]), .Z(n29640)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    LUT4 i15204_2_lut_3_lut (.A(n1294[0]), .B(n1294[8]), .C(\select[7] ), 
         .Z(n15879)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15204_2_lut_3_lut.init = 16'h1010;
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n2036[0]), .SP(n31750), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    LUT4 i15203_2_lut_3_lut (.A(n1294[0]), .B(n1294[8]), .C(\select[2] ), 
         .Z(n15885)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15203_2_lut_3_lut.init = 16'h1010;
    FD1S3IX bufcount__i0 (.D(n15872), .CK(debug_c_c), .CD(n33455), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n30802), .SP(n13568), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    LUT4 esc_data_1__bdd_4_lut (.A(esc_data[1]), .B(esc_data[3]), .C(esc_data[2]), 
         .D(esc_data[4]), .Z(n30672)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)))+!A (B+(C+(D)))) */ ;
    defparam esc_data_1__bdd_4_lut.init = 16'hd7fe;
    LUT4 i1_2_lut_3_lut_adj_61 (.A(n1294[0]), .B(n1294[8]), .C(\select[4] ), 
         .Z(n29639)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_61.init = 16'h1010;
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2619), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i4 (.D(n5604[4]), .SP(n13568), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n5604[2]), .SP(n13568), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n5604[1]), .SP(n13568), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    LUT4 Select_4192_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[6] ), .D(n33446), .Z(n2)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4192_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2617), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i3 (.D(n31887), .CK(debug_c_c), .CD(n33455), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n33438), .CK(debug_c_c), .CD(n33455), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n15046), .CK(debug_c_c), .CD(n33455), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3IX buffer_0___i1 (.D(n28985), .SP(n21320), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 Select_4195_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[3] ), .D(rw), .Z(n2_adj_43)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4195_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX tx_data_i0_i4 (.D(n2036[4]), .SP(n31750), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2036[3]), .SP(n31750), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_62 (.A(register_addr[2]), .B(register_addr[5]), .C(\register[2][0] ), 
         .D(n29956), .Z(n29428)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_62.init = 16'h0010;
    LUT4 i22804_3_lut (.A(register_addr_c[6]), .B(\register_addr[3] ), .C(register_addr_c[7]), 
         .Z(n29956)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22804_3_lut.init = 16'hfefe;
    FD1P3AX tx_data_i0_i1 (.D(n2036[1]), .SP(n31750), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_293_3_lut (.A(\select[4] ), .B(n31765), .C(rw), 
         .Z(n31716)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_293_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_adj_63 (.A(\register_addr[1] ), .B(\steps_reg[5] ), .Z(n14)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_63.init = 16'h8888;
    LUT4 Select_4194_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[4] ), .D(rw), .Z(n2_adj_44)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4194_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut (.A(n31827), .B(n27707), .C(n31720), .D(n33447), 
         .Z(n14124)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut.init = 16'hff20;
    LUT4 Select_4191_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[7] ), .D(rw), .Z(n2_adj_45)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4191_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1S3IX state_FSM_i21 (.D(n11867), .CK(debug_c_c), .CD(n31751), .Q(n1306));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    LUT4 Select_4196_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[2] ), .D(rw), .Z(n2_adj_46)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4196_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1S3IX state_FSM_i20 (.D(n10734), .CK(debug_c_c), .CD(n31751), .Q(n1294[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n29123), .CK(debug_c_c), .CD(n31751), .Q(n1294[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n11865), .CK(debug_c_c), .CD(n31751), .Q(n1309));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n10743), .CK(debug_c_c), .CD(n31751), .Q(n1294[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1406), .CK(debug_c_c), .CD(n31751), .Q(n1294[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1405), .CK(debug_c_c), .CD(n31751), .Q(n1312));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1294[12]), .CK(debug_c_c), .CD(n31751), 
            .Q(n1294[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1294[11]), .CK(debug_c_c), .CD(n31751), 
            .Q(n1294[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1294[10]), .CK(debug_c_c), .CD(n31751), 
            .Q(n1294[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1399), .CK(debug_c_c), .CD(n31751), .Q(n1294[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1294[8]), .CK(debug_c_c), .CD(n31751), 
            .Q(n1294[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1294[7]), .CK(debug_c_c), .CD(n31751), .Q(n1294[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1294[6]), .CK(debug_c_c), .CD(n31751), .Q(n1294[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1294[5]), .CK(debug_c_c), .CD(n31751), .Q(n1294[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n29655), .CK(debug_c_c), .CD(n31751), .Q(n1294[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n29418), .CK(debug_c_c), .CD(n31751), .Q(n1294[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n11698), .CK(debug_c_c), .CD(n31751), .Q(n1294[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n29153), .CK(debug_c_c), .CD(n31751), .Q(n1294[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i2 (.D(n29187), .CK(debug_c_c), .CD(n31751), .Q(n1294[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    LUT4 Select_4197_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[1] ), .D(rw), .Z(n2_adj_47)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4197_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3IX sendcount__i4 (.D(n31236), .SP(n31757), .CD(n31728), .CK(debug_c_c), 
            .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 Select_4198_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[0] ), .D(rw), .Z(n2_adj_48)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4198_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_64 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29708)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_64.init = 16'hfbfb;
    LUT4 Select_4193_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31765), 
         .C(\read_value[5] ), .D(n33446), .Z(n2_adj_49)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4193_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_65 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29709)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_65.init = 16'hbfbf;
    LUT4 i23149_2_lut_rep_275_3_lut_4_lut (.A(rw), .B(n31717), .C(register_addr[0]), 
         .D(n31867), .Z(n31698)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i23149_2_lut_rep_275_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_adj_66 (.A(rx_data[1]), .B(rx_data[4]), .Z(n29632)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_66.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(n31807), .C(n191), 
         .D(\register_addr[1] ), .Z(n29590)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i4415_2_lut_rep_276_3_lut_4_lut (.A(rw), .B(n31717), .C(register_addr[0]), 
         .D(n31867), .Z(n31699)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4415_2_lut_rep_276_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_3_lut_rep_282_4_lut (.A(register_addr[2]), .B(n31807), .C(n31822), 
         .D(n13671), .Z(n31705)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_rep_282_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_3_lut_4_lut_adj_67 (.A(register_addr[2]), .B(n31807), 
         .C(n191), .D(\register_addr[1] ), .Z(n8940)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_67.init = 16'h0010;
    LUT4 i22965_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n31874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22965_then_3_lut.init = 16'hcaca;
    LUT4 i22965_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n31873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22965_else_3_lut.init = 16'hcaca;
    LUT4 i22968_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n31877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22968_then_3_lut.init = 16'hcaca;
    LUT4 i22968_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n31876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22968_else_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(\select[4] ), .B(n31765), .C(prev_select), 
         .D(n33447), .Z(n2658)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_3_lut_4_lut (.A(register_addr[2]), .B(n31807), .C(n21), .D(n31822), 
         .Z(n29452)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_4_lut.init = 16'h0010;
    FD1P3IX sendcount__i3 (.D(n19[3]), .SP(n31757), .CD(n31728), .CK(debug_c_c), 
            .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3IX sendcount__i2 (.D(n19[2]), .SP(n31757), .CD(n31728), .CK(debug_c_c), 
            .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n19[1]), .SP(n31757), .CD(n31728), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_68 (.A(register_addr[0]), .B(n31745), .C(n185), 
         .D(n33447), .Z(n14252)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_68.init = 16'hff10;
    LUT4 i1_2_lut_adj_69 (.A(rx_data[0]), .B(rx_data[5]), .Z(n29623)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_69.init = 16'h2222;
    LUT4 i15_2_lut_rep_323_4_lut (.A(n31806), .B(\register_addr[4] ), .C(select[3]), 
         .D(rw), .Z(n31746)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i15_2_lut_rep_323_4_lut.init = 16'h4000;
    LUT4 i22971_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n31880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22971_then_3_lut.init = 16'hcaca;
    LUT4 i22971_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n31879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22971_else_3_lut.init = 16'hcaca;
    LUT4 i23218_4_lut (.A(debug_c_7), .B(n29623), .C(n1294[3]), .D(n4_c), 
         .Z(n29418)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i23218_4_lut.init = 16'h20a0;
    LUT4 i1_2_lut_4_lut_adj_70 (.A(prev_select), .B(n31723), .C(n29710), 
         .D(n33447), .Z(n13757)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_70.init = 16'hff04;
    LUT4 i1_2_lut_4_lut_adj_71 (.A(n31779), .B(n13671), .C(n31822), .D(\register_addr[1] ), 
         .Z(n29552)) /* synthesis lut_function=(!(A (B+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_71.init = 16'h3700;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n31883)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i1_4_lut (.A(escape), .B(rx_data[7]), .C(rx_data[6]), .D(n31238), 
         .Z(n4_c)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n31882)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 i5296_3_lut (.A(debug_c_7), .B(n1294[3]), .C(n1294[2]), .Z(n11698)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5296_3_lut.init = 16'h5454;
    LUT4 i8638_then_4_lut (.A(bufcount[3]), .B(n1294[0]), .C(n1294[3]), 
         .D(n1294[4]), .Z(n31886)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8638_then_4_lut.init = 16'haaa2;
    LUT4 i8638_else_4_lut (.A(bufcount[3]), .B(n1294[0]), .C(n1294[3]), 
         .D(n1294[4]), .Z(n31885)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8638_else_4_lut.init = 16'h0002;
    LUT4 i23399_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n31889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23399_then_3_lut.init = 16'hcaca;
    LUT4 i23399_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n31888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23399_else_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_72 (.A(n1294[4]), .B(debug_c_7), .C(n1294[2]), .D(n29419), 
         .Z(n29153)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_72.init = 16'heeea;
    LUT4 i1_4_lut_adj_73 (.A(n15), .B(n1294[3]), .C(n1294[0]), .D(n30012), 
         .Z(n29419)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_73.init = 16'h50dc;
    LUT4 i22860_3_lut (.A(n13070), .B(escape), .C(n15), .Z(n30012)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i22860_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_3_lut_adj_74 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29758)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_74.init = 16'hfbfb;
    LUT4 i22884_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n31892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22884_then_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_75 (.A(n31795), .B(debug_c_7), .C(n13182), .D(n8), 
         .Z(n29187)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_75.init = 16'hdc50;
    LUT4 i22884_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n31891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22884_else_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(n15), .B(n1294[1]), .C(n1294[0]), .Z(n8)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i22956_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n31901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22956_then_3_lut.init = 16'hcaca;
    LUT4 i22956_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n31900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22956_else_3_lut.init = 16'hcaca;
    LUT4 i15_2_lut_3_lut_4_lut (.A(\register_addr[4] ), .B(n31806), .C(rw), 
         .D(select[3]), .Z(n47)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;
    defparam i15_2_lut_3_lut_4_lut.init = 16'hd000;
    LUT4 Select_4201_i6_2_lut_3_lut_4_lut (.A(\register_addr[4] ), .B(n31806), 
         .C(\read_size[2] ), .D(select[3]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;
    defparam Select_4201_i6_2_lut_3_lut_4_lut.init = 16'hd000;
    LUT4 Select_4197_i4_2_lut_3_lut_4_lut (.A(n31739), .B(\select[4] ), 
         .C(\read_value[1]_adj_50 ), .D(rw), .Z(n4)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_4197_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i22959_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n31904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22959_then_3_lut.init = 16'hcaca;
    LUT4 i22959_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n31903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22959_else_3_lut.init = 16'hcaca;
    LUT4 n30016_bdd_4_lut (.A(bufcount[1]), .B(n1294[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n32225)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n30016_bdd_4_lut.init = 16'h0080;
    LUT4 i2_3_lut_4_lut_adj_76 (.A(n31739), .B(\select[4] ), .C(n27707), 
         .D(n29699), .Z(n3970)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_76.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_77 (.A(register_addr[5]), .B(n31807), 
         .C(\register_addr[1] ), .D(n160), .Z(n78)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_77.init = 16'h0100;
    LUT4 i2_3_lut_rep_340_4_lut (.A(register_addr[5]), .B(n31807), .C(register_addr[2]), 
         .D(\select[4] ), .Z(n31763)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_340_4_lut.init = 16'h0100;
    FD1S3AX escape_501 (.D(n10514), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_78 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29757)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_78.init = 16'hbfbf;
    LUT4 Select_4157_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[19] ), .Z(n3)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4157_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 Select_4154_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[20] ), .Z(n3_adj_51)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4154_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_79 (.A(register_addr[5]), .B(n31807), 
         .C(\read_size[2]_adj_52 ), .D(n160), .Z(n20)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_79.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_80 (.A(register_addr[5]), .B(n31807), .C(n31832), 
         .D(register_addr[2]), .Z(n29808)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_80.init = 16'h1110;
    LUT4 i1_2_lut_rep_316_3_lut_4_lut (.A(register_addr[5]), .B(n31807), 
         .C(register_addr[2]), .D(\register_addr[4] ), .Z(n31739)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_316_3_lut_4_lut.init = 16'hfffe;
    LUT4 i14798_4_lut (.A(sendcount[3]), .B(n9_adj_74), .C(sendcount[2]), 
         .D(n31830), .Z(n19[3])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(271[10:37])
    defparam i14798_4_lut.init = 16'h4888;
    LUT4 Select_4151_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[21] ), .Z(n3_adj_53)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4151_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_81 (.A(n1294[16]), .B(n1294[19]), .Z(n2045)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_81.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_82 (.A(n31827), .B(prev_select_adj_54), .C(n31706), 
         .D(n33447), .Z(n14172)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_82.init = 16'hff02;
    LUT4 Select_4148_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[22] ), .Z(n3_adj_55)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4148_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 Select_4145_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[23] ), .Z(n3_adj_56)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4145_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 Select_4142_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[24] ), .Z(n3_adj_57)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4142_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 Select_4139_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[25] ), .Z(n3_adj_58)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4139_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_83 (.A(n1294[4]), .B(\buffer[0] [1]), .C(n11_adj_81), 
         .D(n14_adj_82), .Z(n28977)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_83.init = 16'heca0;
    LUT4 n12791_bdd_2_lut_23502 (.A(sendcount[0]), .B(sendcount[3]), .Z(n30796)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n12791_bdd_2_lut_23502.init = 16'hbbbb;
    FD1P3AX rw_498 (.D(n1294[10]), .SP(n2617), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_84 (.A(n1294[4]), .B(\buffer[0] [2]), .C(n11_adj_83), 
         .D(n14_adj_82), .Z(n28981)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_84.init = 16'heca0;
    LUT4 Select_4136_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[26] ), .Z(n3_adj_59)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4136_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_85 (.A(n1294[4]), .B(\buffer[0] [3]), .C(n11_adj_85), 
         .D(n14_adj_82), .Z(n28983)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_85.init = 16'heca0;
    LUT4 Select_4133_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[27] ), .Z(n3_adj_60)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4133_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_86 (.A(n1294[4]), .B(\buffer[0] [4]), .C(n11_adj_87), 
         .D(n14_adj_82), .Z(n28991)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_86.init = 16'heca0;
    LUT4 Select_4130_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[28] ), .Z(n3_adj_61)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4130_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 n32223_bdd_4_lut (.A(n32223), .B(n1294[4]), .C(n32225), .D(bufcount[2]), 
         .Z(n33438)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n32223_bdd_4_lut.init = 16'heef0;
    LUT4 i1_4_lut_adj_87 (.A(n1294[4]), .B(\buffer[0] [5]), .C(n11_adj_89), 
         .D(n14_adj_82), .Z(n28989)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_87.init = 16'heca0;
    LUT4 Select_4127_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[29] ), .Z(n3_adj_62)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4127_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_88 (.A(n1294[4]), .B(\buffer[0] [6]), .C(n11_adj_91), 
         .D(n14_adj_82), .Z(n28987)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_88.init = 16'heca0;
    LUT4 i1_4_lut_adj_89 (.A(n1294[4]), .B(\buffer[0] [7]), .C(n11_adj_92), 
         .D(n14_adj_82), .Z(n29059)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_89.init = 16'heca0;
    LUT4 Select_4124_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[30] ), .Z(n3_adj_63)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4124_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_rep_342_4_lut (.A(register_addr[5]), .B(n31807), .C(register_addr[2]), 
         .D(\register_addr[4] ), .Z(n31765)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_342_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_318_3_lut_4_lut (.A(register_addr[5]), .B(n31807), 
         .C(\select[4] ), .D(n160), .Z(n31741)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_318_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4121_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[31] ), .Z(n3_adj_64)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4121_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 Select_4160_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[18] ), .Z(n3_adj_65)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4160_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_90 (.A(n1294[4]), .B(\buffer[1] [0]), .C(n11_adj_96), 
         .D(n14_adj_82), .Z(n28979)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_90.init = 16'heca0;
    LUT4 Select_4163_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[17] ), .Z(n3_adj_66)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4163_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_91 (.A(n31815), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n13182), .Z(n29655)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_91.init = 16'h0e00;
    LUT4 Select_4166_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[16] ), .Z(n3_adj_67)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4166_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n31815), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_adj_99)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_92 (.A(bufcount[0]), .B(n31815), .C(\buffer[0] [1]), 
         .D(rx_data[1]), .Z(n11_adj_81)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_92.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_93 (.A(bufcount[0]), .B(n31815), .C(\buffer[0] [2]), 
         .D(rx_data[2]), .Z(n11_adj_83)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_93.init = 16'hf1e0;
    LUT4 Select_4169_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[15] ), .Z(n3_adj_68)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4169_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i24_3_lut_4_lut_adj_94 (.A(bufcount[0]), .B(n31815), .C(\buffer[0] [3]), 
         .D(rx_data[3]), .Z(n11_adj_85)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_94.init = 16'hf1e0;
    LUT4 Select_4172_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[14] ), .Z(n3_adj_69)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4172_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i24_3_lut_4_lut_adj_95 (.A(bufcount[0]), .B(n31815), .C(rx_data[4]), 
         .D(\buffer[0] [4]), .Z(n11_adj_87)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_95.init = 16'hfe10;
    LUT4 i1_4_lut_adj_96 (.A(n1294[4]), .B(\buffer[1] [1]), .C(n11_adj_102), 
         .D(n14_adj_82), .Z(n28959)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_96.init = 16'heca0;
    LUT4 i9211_4_lut (.A(escape), .B(n13070), .C(n6_adj_103), .D(n1294[3]), 
         .Z(n10514)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i9211_4_lut.init = 16'h1aaa;
    LUT4 i1_4_lut_adj_97 (.A(n1294[4]), .B(\buffer[1] [2]), .C(n11_adj_104), 
         .D(n14_adj_82), .Z(n29039)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_97.init = 16'heca0;
    LUT4 Select_4175_i3_2_lut_4_lut (.A(n31754), .B(rw), .C(\select[4] ), 
         .D(\read_value[13] ), .Z(n3_adj_70)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4175_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i24_3_lut_4_lut_adj_98 (.A(bufcount[0]), .B(n31815), .C(rx_data[5]), 
         .D(\buffer[0] [5]), .Z(n11_adj_89)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_98.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_99 (.A(bufcount[0]), .B(n31815), .C(\buffer[0] [6]), 
         .D(rx_data[6]), .Z(n11_adj_91)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_99.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_100 (.A(n1294[4]), .B(\buffer[1] [3]), .C(n11_adj_106), 
         .D(n14_adj_82), .Z(n29055)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_100.init = 16'heca0;
    LUT4 i2_2_lut (.A(debug_c_7), .B(n31783), .Z(n6_adj_103)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i24_3_lut_4_lut_adj_101 (.A(bufcount[0]), .B(n31815), .C(rx_data[7]), 
         .D(\buffer[0] [7]), .Z(n11_adj_92)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_101.init = 16'hfe10;
    LUT4 i1_4_lut_adj_102 (.A(n1294[4]), .B(\buffer[1] [4]), .C(n11_adj_107), 
         .D(n14_adj_82), .Z(n29095)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_102.init = 16'heca0;
    LUT4 i1_4_lut_adj_103 (.A(n1294[4]), .B(\buffer[1] [5]), .C(n11_adj_108), 
         .D(n14_adj_82), .Z(n29047)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_103.init = 16'heca0;
    LUT4 i1_4_lut_adj_104 (.A(n1294[4]), .B(\buffer[1] [6]), .C(n11_adj_109), 
         .D(n14_adj_82), .Z(n29011)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_104.init = 16'heca0;
    LUT4 i1_4_lut_adj_105 (.A(n1294[4]), .B(\buffer[1] [7]), .C(n11_adj_110), 
         .D(n14_adj_82), .Z(n28969)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_105.init = 16'heca0;
    LUT4 i2_4_lut (.A(databus[0]), .B(n5), .C(n1294[13]), .D(n29523), 
         .Z(n28079)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 select_2068_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1294[4]), 
         .C(rx_data[0]), .D(n29758), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n31829), .B(n31805), .C(n4_adj_111), 
         .D(n31893), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i2_4_lut_adj_106 (.A(databus[1]), .B(n5_adj_112), .C(n1294[13]), 
         .D(n29532), .Z(n28074)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_106.init = 16'hffec;
    LUT4 select_2068_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1294[4]), 
         .C(rx_data[1]), .D(n29758), .Z(n5_adj_112)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_107 (.A(databus[2]), .B(n5_adj_113), .C(n1294[13]), 
         .D(n29522), .Z(n28077)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_107.init = 16'hffec;
    LUT4 Select_4178_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[12] ), .Z(n3_adj_71)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4178_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 select_2068_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1294[4]), 
         .C(rx_data[2]), .D(n29758), .Z(n5_adj_113)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4181_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[11] ), .Z(n3_adj_72)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4181_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n31829), .B(n31805), .C(n4_adj_116), 
         .D(n31881), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 Select_4184_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[10] ), .Z(n3_adj_73)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4184_i3_2_lut_4_lut.init = 16'h8000;
    FD1P3IX send_491 (.D(n33445), .SP(n2045), .CD(n28025), .CK(debug_c_c), 
            .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n31829), .B(n31805), .C(n4_adj_118), 
         .D(n31875), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_rep_462 (.A(\register_addr[4] ), .B(n31787), .C(n31828), 
         .D(register_addr[2]), .Z(n33457)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_462.init = 16'hffef;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1294[4]), .B(n31817), .C(bufcount[0]), 
         .D(n31781), .Z(n28097)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hd222;
    LUT4 n30800_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n31834), .C(n31890), 
         .D(n30800), .Z(n30801)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n30800_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 i22962_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n31871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22962_then_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n31829), .B(n31805), .C(n4_adj_119), 
         .D(n31902), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n31829), .B(n31805), .C(n4_adj_120), 
         .D(n31905), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n31829), .B(n31805), .C(n4_adj_121), 
         .D(n31872), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n31829), .B(n31805), .C(n4_adj_122), 
         .D(n31878), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i2_3_lut (.A(n15_adj_123), .B(register_addr[0]), .C(\register_addr[4] ), 
         .Z(n28937)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i2_3_lut.init = 16'h0202;
    LUT4 i2_3_lut_rep_357_4_lut (.A(register_addr[5]), .B(n31840), .C(select[3]), 
         .D(\register_addr[4] ), .Z(n31780)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_rep_357_4_lut.init = 16'h1000;
    LUT4 i2_4_lut_adj_108 (.A(databus[3]), .B(n5_adj_124), .C(n1294[13]), 
         .D(n29524), .Z(n28075)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_108.init = 16'hffec;
    LUT4 Select_4187_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[9] ), .Z(n3_adj_74)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4187_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i20566_2_lut (.A(n33446), .B(prev_select_adj_54), .Z(n27707)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20566_2_lut.init = 16'heeee;
    LUT4 i23146_2_lut_3_lut_4_lut (.A(n31867), .B(n31706), .C(n33447), 
         .D(register_addr[0]), .Z(n22093)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam i23146_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 Select_4190_i3_2_lut_4_lut (.A(n31754), .B(n33446), .C(\select[4] ), 
         .D(\read_value[8] ), .Z(n3_adj_75)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4190_i3_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_339_3_lut_4_lut (.A(register_addr[5]), .B(n31840), 
         .C(select[3]), .D(\register_addr[4] ), .Z(n31762)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i1_2_lut_rep_339_3_lut_4_lut.init = 16'he0f0;
    LUT4 select_2068_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1294[4]), 
         .C(rx_data[3]), .D(n29758), .Z(n5_adj_124)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_109 (.A(databus[4]), .B(n5_adj_127), .C(n1294[13]), 
         .D(n29525), .Z(n28076)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_109.init = 16'hffec;
    LUT4 select_2068_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1294[4]), 
         .C(rx_data[4]), .D(n29758), .Z(n5_adj_127)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_322_3_lut_4_lut (.A(\register_addr[3] ), .B(n31840), 
         .C(\register_addr[1] ), .D(register_addr[2]), .Z(n31745)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_322_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_110 (.A(databus[5]), .B(n5_adj_128), .C(n1294[13]), 
         .D(n29526), .Z(n28072)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_110.init = 16'hffec;
    LUT4 select_2068_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1294[4]), 
         .C(rx_data[5]), .D(n29758), .Z(n5_adj_128)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_331_3_lut_4_lut (.A(\register_addr[3] ), .B(n31840), 
         .C(n160), .D(register_addr[5]), .Z(n31754)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_331_3_lut_4_lut.init = 16'h0010;
    LUT4 i22678_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n31739), .C(prev_select_adj_76), 
         .D(register_addr[0]), .Z(n29823)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22678_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_111 (.A(databus[6]), .B(n5_adj_130), .C(n1294[13]), 
         .D(n29527), .Z(n28091)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_111.init = 16'hffec;
    LUT4 i1_2_lut_rep_280_3_lut_4_lut (.A(register_addr[2]), .B(n31772), 
         .C(n33446), .D(\select[4] ), .Z(n31703)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_280_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_349_3_lut_4_lut (.A(\register_addr[3] ), .B(n31840), 
         .C(\register_addr[4] ), .D(register_addr[5]), .Z(n31772)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_349_3_lut_4_lut.init = 16'hfffe;
    LUT4 select_2068_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1294[4]), 
         .C(rx_data[6]), .D(n29758), .Z(n5_adj_130)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_295_4_lut (.A(register_addr[2]), .B(n31772), .C(register_addr[0]), 
         .D(\register_addr[1] ), .Z(n31718)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_295_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_351_3_lut_4_lut (.A(\register_addr[3] ), .B(n31840), 
         .C(n160), .D(register_addr[5]), .Z(n31774)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_351_3_lut_4_lut.init = 16'h1000;
    LUT4 i9640_4_lut_4_lut (.A(\register_addr[1] ), .B(n31739), .C(register_addr[0]), 
         .D(n14022), .Z(n16046)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+(C+!(D))))) */ ;
    defparam i9640_4_lut_4_lut.init = 16'h2300;
    LUT4 i2_4_lut_adj_112 (.A(databus[7]), .B(n5_adj_131), .C(n1294[13]), 
         .D(n29528), .Z(n28073)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_112.init = 16'hffec;
    LUT4 select_2068_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1294[4]), 
         .C(rx_data[7]), .D(n29758), .Z(n5_adj_131)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 i9639_3_lut_4_lut (.A(register_addr[2]), .B(n31772), .C(n31828), 
         .D(n14022), .Z(n16045)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i9639_3_lut_4_lut.init = 16'hfe00;
    LUT4 i2_4_lut_adj_113 (.A(databus[8]), .B(n5_adj_132), .C(n1294[13]), 
         .D(n29529), .Z(n28034)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_113.init = 16'hffec;
    LUT4 select_2068_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1294[4]), 
         .C(rx_data[0]), .D(n29757), .Z(n5_adj_132)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 n29626_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n30673)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n29626_bdd_4_lut.init = 16'h4001;
    LUT4 i23168_3_lut_4_lut (.A(n12_c), .B(\buffer[0] [2]), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n29767)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23168_3_lut_4_lut.init = 16'h4000;
    LUT4 i23205_3_lut_4_lut (.A(n12_c), .B(\buffer[0] [2]), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n29766)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23205_3_lut_4_lut.init = 16'h0004;
    LUT4 i23189_3_lut_4_lut (.A(\buffer[0] [2]), .B(n12_c), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n28151)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23189_3_lut_4_lut.init = 16'h0010;
    LUT4 \buffer_0[[1__bdd_4_lut_23743  (.A(\buffer[0] [1]), .B(n29744), 
         .C(n29640), .D(n1747), .Z(n31686)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam \buffer_0[[1__bdd_4_lut_23743 .init = 16'h22f0;
    LUT4 i2_1_lut_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(n31772), .C(register_addr[0]), 
         .D(\register_addr[1] ), .Z(n24748)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i2_1_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_114 (.A(register_addr[2]), .B(n31772), 
         .C(register_addr[0]), .D(\register_addr[1] ), .Z(n250)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_114.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_115 (.A(\buffer[0] [2]), .B(n12_c), .C(\buffer[0] [0]), 
         .Z(n29744)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i1_2_lut_3_lut_adj_115.init = 16'hefef;
    LUT4 \buffer_0[[1__bdd_4_lut  (.A(\buffer[0] [1]), .B(n29744), .C(n15875), 
         .D(n1747), .Z(n31687)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam \buffer_0[[1__bdd_4_lut .init = 16'h11f0;
    LUT4 i1_2_lut_adj_116 (.A(\register_addr[4] ), .B(register_addr[2]), 
         .Z(n160)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_116.init = 16'h2222;
    LUT4 i2_4_lut_adj_117 (.A(databus[9]), .B(n5_adj_133), .C(n1294[13]), 
         .D(n29531), .Z(n28086)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_117.init = 16'hffec;
    LUT4 select_2068_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1294[4]), 
         .C(rx_data[1]), .D(n29757), .Z(n5_adj_133)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_118 (.A(databus[10]), .B(n5_adj_134), .C(n1294[13]), 
         .D(n29521), .Z(n27895)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_118.init = 16'hffec;
    LUT4 select_2068_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1294[4]), 
         .C(rx_data[2]), .D(n29757), .Z(n5_adj_134)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i24_3_lut_4_lut_adj_119 (.A(bufcount[0]), .B(n31815), .C(\buffer[1] [0]), 
         .D(rx_data[0]), .Z(n11_adj_96)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_119.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_120 (.A(bufcount[0]), .B(n31815), .C(\buffer[1] [1]), 
         .D(rx_data[1]), .Z(n11_adj_102)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_120.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_121 (.A(bufcount[0]), .B(n31815), .C(\buffer[1] [2]), 
         .D(rx_data[2]), .Z(n11_adj_104)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_121.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_122 (.A(bufcount[0]), .B(n31815), .C(rx_data[3]), 
         .D(\buffer[1] [3]), .Z(n11_adj_106)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_122.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_123 (.A(bufcount[0]), .B(n31815), .C(rx_data[4]), 
         .D(\buffer[1] [4]), .Z(n11_adj_107)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_123.init = 16'hfd20;
    LUT4 i2_4_lut_adj_124 (.A(databus[11]), .B(n5_adj_135), .C(n1294[13]), 
         .D(n29516), .Z(n28005)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_124.init = 16'hffec;
    LUT4 select_2068_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1294[4]), 
         .C(rx_data[3]), .D(n29757), .Z(n5_adj_135)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i22787_2_lut_rep_283_3_lut_4_lut (.A(register_addr[2]), .B(n31772), 
         .C(rw), .D(\register_addr[1] ), .Z(n31706)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22787_2_lut_rep_283_3_lut_4_lut.init = 16'hfffe;
    LUT4 i24_3_lut_4_lut_adj_125 (.A(bufcount[0]), .B(n31815), .C(rx_data[5]), 
         .D(\buffer[1] [5]), .Z(n11_adj_108)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_125.init = 16'hfd20;
    LUT4 i2_4_lut_adj_126 (.A(databus[12]), .B(n5_adj_136), .C(n1294[13]), 
         .D(n29534), .Z(n28083)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_126.init = 16'hffec;
    LUT4 i24_3_lut_4_lut_adj_127 (.A(bufcount[0]), .B(n31815), .C(\buffer[1] [6]), 
         .D(rx_data[6]), .Z(n11_adj_109)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_127.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_128 (.A(bufcount[0]), .B(n31815), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_110)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_128.init = 16'hf2d0;
    LUT4 select_2068_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1294[4]), 
         .C(rx_data[4]), .D(n29757), .Z(n5_adj_136)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 i22962_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n31870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22962_else_3_lut.init = 16'hcaca;
    LUT4 i3190_2_lut_rep_392 (.A(bufcount[1]), .B(bufcount[2]), .Z(n31815)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3190_2_lut_rep_392.init = 16'heeee;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n31750), .CD(n16067), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    LUT4 i2824_2_lut_rep_372_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n31795)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2824_2_lut_rep_372_3_lut.init = 16'hfefe;
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n31750), .CD(n16067), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    LUT4 i902_2_lut_rep_393 (.A(escape), .B(debug_c_7), .Z(n31816)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i902_2_lut_rep_393.init = 16'hbbbb;
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n31750), .CD(n16067), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_358_4_lut (.A(escape), .B(debug_c_7), .C(n30016), 
         .D(n1294[4]), .Z(n31781)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_358_4_lut.init = 16'hfffb;
    LUT4 i2_4_lut_adj_129 (.A(databus[13]), .B(n5_adj_137), .C(n1294[13]), 
         .D(n29530), .Z(n28022)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_129.init = 16'hffec;
    LUT4 i15554_3_lut_rep_394 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n31817)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15554_3_lut_rep_394.init = 16'hecec;
    LUT4 i2_2_lut_rep_381_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1294[4]), .Z(n31804)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_381_4_lut.init = 16'hecff;
    LUT4 sendcount_1__bdd_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(sendcount[3]), 
         .D(sendcount[2]), .Z(n31235)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_1__bdd_4_lut.init = 16'h6aaa;
    LUT4 i1_2_lut_4_lut_adj_130 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1294[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_130.init = 16'hec00;
    LUT4 select_2068_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1294[4]), 
         .C(rx_data[5]), .D(n29757), .Z(n5_adj_137)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4197_i1_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31774), 
         .C(\read_value[1]_adj_77 ), .D(rw), .Z(n1)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4197_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 sendcount_4__bdd_3_lut (.A(sendcount[4]), .B(n31235), .C(\sendcount[1] ), 
         .Z(n31236)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut.init = 16'hcaca;
    LUT4 rx_data_2__bdd_4_lut (.A(rx_data[2]), .B(rx_data[3]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n31238)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_2__bdd_4_lut.init = 16'h6001;
    LUT4 i2_4_lut_adj_131 (.A(databus[14]), .B(n5_adj_139), .C(n1294[13]), 
         .D(n29519), .Z(n28008)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_131.init = 16'hffec;
    LUT4 select_2068_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1294[4]), 
         .C(rx_data[6]), .D(n29757), .Z(n5_adj_139)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_132 (.A(databus[15]), .B(n5_adj_140), .C(n1294[13]), 
         .D(n29536), .Z(n28084)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_132.init = 16'hffec;
    LUT4 select_2068_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1294[4]), 
         .C(rx_data[7]), .D(n29757), .Z(n5_adj_140)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_399 (.A(\register_addr[4] ), .B(register_addr[5]), 
         .Z(n31822)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_399.init = 16'heeee;
    LUT4 i2_4_lut_adj_133 (.A(databus[16]), .B(n5_adj_141), .C(n1294[13]), 
         .D(n29535), .Z(n28082)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_133.init = 16'hffec;
    LUT4 select_2068_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1294[4]), 
         .C(rx_data[0]), .D(n29708), .Z(n5_adj_141)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_134 (.A(\register_addr[4] ), .B(register_addr[5]), 
         .C(n31840), .D(\register_addr[3] ), .Z(n29738)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_134.init = 16'hfffe;
    LUT4 i15521_3_lut_rep_327 (.A(n2557), .B(n31783), .C(n1294[18]), .Z(n31750)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15521_3_lut_rep_327.init = 16'hc8c8;
    LUT4 i4_2_lut_rep_400 (.A(n1312), .B(n1294[15]), .Z(n31823)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_400.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_135 (.A(n1312), .B(n1294[15]), .C(n1294[12]), 
         .Z(n29795)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_135.init = 16'hfefe;
    LUT4 i1_2_lut_rep_401 (.A(n1294[3]), .B(n1294[19]), .Z(n31824)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_401.init = 16'heeee;
    LUT4 i23100_2_lut_3_lut (.A(n2557), .B(n31783), .C(n1294[18]), .Z(n16067)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i23100_2_lut_3_lut.init = 16'h0808;
    PFUMX i8640 (.BLUT(n15045), .ALUT(n1690[1]), .C0(n1695), .Z(n15046));
    LUT4 i1_2_lut_rep_402 (.A(n1294[11]), .B(n1294[9]), .Z(n31825)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_402.init = 16'heeee;
    LUT4 i3_2_lut_3_lut_4_lut (.A(n1294[11]), .B(n1294[9]), .C(n1294[19]), 
         .D(n1294[3]), .Z(n9_adj_142)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_4_lut (.A(n1294[7]), .B(n1294[13]), .C(n1294[5]), .D(n1309), 
         .Z(n8_adj_143)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut_4_lut.init = 16'hfffe;
    PFUMX i9466 (.BLUT(n15871), .ALUT(n28097), .C0(n1695), .Z(n15872));
    LUT4 i1_2_lut_4_lut_adj_136 (.A(n1294[7]), .B(n1294[13]), .C(n1294[5]), 
         .D(n1294[6]), .Z(n6_adj_144)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_4_lut_adj_136.init = 16'hfffe;
    LUT4 i1_2_lut_adj_137 (.A(\register_addr[4] ), .B(register_addr[5]), 
         .Z(n191)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_137.init = 16'h8888;
    LUT4 i2_4_lut_adj_138 (.A(databus[17]), .B(n5_adj_145), .C(n1294[13]), 
         .D(n29533), .Z(n28048)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_138.init = 16'hffec;
    LUT4 i1_2_lut_adj_139 (.A(\register_addr[1] ), .B(\steps_reg[6] ), .Z(n13)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_139.init = 16'h8888;
    LUT4 i1_2_lut_rep_403 (.A(\register_addr[1] ), .B(\select[4] ), .Z(n31826)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_403.init = 16'h8888;
    LUT4 i2_3_lut_rep_301_4_lut (.A(\register_addr[1] ), .B(\select[4] ), 
         .C(n29874), .D(\register_addr[4] ), .Z(n31724)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_301_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_rep_404 (.A(register_addr[0]), .B(\select[4] ), .Z(n31827)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_404.init = 16'h4444;
    LUT4 select_2068_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1294[4]), 
         .C(rx_data[1]), .D(n29708), .Z(n5_adj_145)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_140 (.A(sendcount[4]), .B(n1_adj_147), .C(n6_adj_148), 
         .D(n12795), .Z(n9_adj_74)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_140.init = 16'hfeff;
    LUT4 i2_3_lut_4_lut_adj_141 (.A(register_addr[0]), .B(\select[4] ), 
         .C(\register_addr[1] ), .D(rw), .Z(n29404)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_141.init = 16'h0004;
    LUT4 i1_2_lut_rep_405 (.A(register_addr[0]), .B(\register_addr[1] ), 
         .Z(n31828)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_405.init = 16'h2222;
    LUT4 equal_52_i1_4_lut (.A(sendcount[0]), .B(n9), .C(n14_adj_78), 
         .D(n10), .Z(n1_adj_147)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_52_i1_4_lut.init = 16'h5556;
    LUT4 i2_4_lut_adj_142 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n31841), .Z(n6_adj_148)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_142.init = 16'he7de;
    LUT4 i23160_2_lut_2_lut_3_lut_4_lut_4_lut_2_lut (.A(\register_addr[1] ), 
         .B(n31739), .Z(n106)) /* synthesis lut_function=(!(A+(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i23160_2_lut_2_lut_3_lut_4_lut_4_lut_2_lut.init = 16'h1111;
    LUT4 i3284_2_lut_rep_406 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n31829)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i3284_2_lut_rep_406.init = 16'h9999;
    LUT4 i14800_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_adj_74), .Z(n19[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i14800_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 n12791_bdd_4_lut_23506_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n30800)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n12791_bdd_4_lut_23506_4_lut.init = 16'h6420;
    LUT4 i1_2_lut_adj_143 (.A(register_addr[0]), .B(\control_reg[7] ), .Z(n8243)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_143.init = 16'h4444;
    LUT4 i3523_2_lut_rep_407 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n31830)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3523_2_lut_rep_407.init = 16'h8888;
    LUT4 i14799_3_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(n9_adj_74), 
         .D(sendcount[2]), .Z(n19[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;
    defparam i14799_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i2_4_lut_adj_144 (.A(databus[18]), .B(n5_adj_151), .C(n1294[13]), 
         .D(n29537), .Z(n28035)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_144.init = 16'hffec;
    LUT4 i54_4_lut (.A(n31739), .B(\read_size[0] ), .C(\read_size[0]_adj_79 ), 
         .D(n31774), .Z(n55)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i54_4_lut.init = 16'hdc50;
    LUT4 select_2068_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1294[4]), 
         .C(rx_data[2]), .D(n29708), .Z(n5_adj_151)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_34_i5_4_lut.init = 16'h88c0;
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2617), .CK(debug_c_c), 
            .Q(register_addr_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2617), .CK(debug_c_c), 
            .Q(register_addr_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2617), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2617), .CK(debug_c_c), 
            .Q(\register_addr[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2617), .CK(debug_c_c), 
            .Q(\register_addr[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2617), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2617), .CK(debug_c_c), 
            .Q(\register_addr[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_145 (.A(\select[4] ), .B(n31739), .C(n20), .D(\read_size[2]_adj_80 ), 
         .Z(n9_adj_81)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_4_lut_adj_145.init = 16'ha2a0;
    LUT4 i2_4_lut_adj_146 (.A(databus[19]), .B(n5_adj_155), .C(n1294[13]), 
         .D(n29538), .Z(n28002)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_146.init = 16'hffec;
    LUT4 i1_2_lut_adj_147 (.A(register_addr[0]), .B(\control_reg[7]_adj_82 ), 
         .Z(n1_adj_83)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_147.init = 16'h4444;
    LUT4 select_2068_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1294[4]), 
         .C(rx_data[3]), .D(n29708), .Z(n5_adj_155)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_35_i5_4_lut.init = 16'h88c0;
    FD1P3IX buffer_0___i2 (.D(n28977), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_148 (.A(databus[20]), .B(n5_adj_158), .C(n1294[13]), 
         .D(n29539), .Z(n28016)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_148.init = 16'hffec;
    LUT4 i3240_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n31781), .C(n31804), 
         .D(bufcount[0]), .Z(n1690[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3240_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    FD1P3IX buffer_0___i3 (.D(n28981), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n28983), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n28991), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n28989), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n28987), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n29059), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n28979), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n28959), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n29039), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n29055), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n29095), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n29047), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n29011), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n28969), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n28079), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n28074), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n28077), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n28075), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n28076), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i22 (.D(n28072), .SP(n9017), .CD(n31751), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    FD1P3IX buffer_0___i23 (.D(n28091), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n28073), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n28034), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n28086), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n27895), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n28005), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n28083), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n28022), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n28008), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n28084), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n28082), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n28048), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n28035), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n28002), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n28016), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n27964), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n28012), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n28030), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n27994), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n27999), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n28013), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n28023), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n28026), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n27998), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n28020), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n28019), .SP(n9017), .CD(n33455), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 select_2068_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1294[4]), 
         .C(rx_data[4]), .D(n29708), .Z(n5_adj_158)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_149 (.A(databus[21]), .B(n5_adj_159), .C(n1294[13]), 
         .D(n29540), .Z(n27964)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_149.init = 16'hffec;
    LUT4 select_2068_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1294[4]), 
         .C(rx_data[5]), .D(n29708), .Z(n5_adj_159)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_150 (.A(databus[22]), .B(n5_adj_160), .C(n1294[13]), 
         .D(n29541), .Z(n28012)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_150.init = 16'hffec;
    LUT4 select_2068_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1294[4]), 
         .C(rx_data[6]), .D(n29708), .Z(n5_adj_160)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_151 (.A(databus[23]), .B(n5_adj_161), .C(n1294[13]), 
         .D(n29542), .Z(n28030)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_151.init = 16'hffec;
    LUT4 select_2068_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1294[4]), 
         .C(rx_data[7]), .D(n29708), .Z(n5_adj_161)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_410 (.A(n1312), .B(sendcount[4]), .Z(n31833)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_410.init = 16'h2222;
    LUT4 motor_pwm_r_c_bdd_2_lut_23346_3_lut (.A(n1312), .B(sendcount[4]), 
         .C(n30673), .Z(n30674)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam motor_pwm_r_c_bdd_2_lut_23346_3_lut.init = 16'h2020;
    PFUMX i23401 (.BLUT(n30801), .ALUT(n30796), .C0(n5613), .Z(n30802));
    LUT4 i14688_2_lut_rep_411 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n31834)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14688_2_lut_rep_411.init = 16'heeee;
    LUT4 i1_2_lut_rep_382_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n31805)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_382_3_lut.init = 16'h1e1e;
    LUT4 i2_4_lut_adj_152 (.A(databus[24]), .B(n5_adj_162), .C(n1294[13]), 
         .D(n29543), .Z(n27994)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_152.init = 16'hffec;
    LUT4 i1_4_lut_adj_153 (.A(n5613), .B(n17[0]), .C(n31783), .D(n1312), 
         .Z(n16049)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_153.init = 16'h8000;
    LUT4 select_2068_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1294[4]), 
         .C(rx_data[0]), .D(n29709), .Z(n5_adj_162)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_122)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_121)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 reduce_or_449_i1_3_lut_4_lut (.A(n31795), .B(n13182), .C(\buffer[0] [7]), 
         .D(n1294[9]), .Z(n1399)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_449_i1_3_lut_4_lut.init = 16'hff80;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_120)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    PFUMX i9474 (.BLUT(n15879), .ALUT(n29767), .C0(n1747), .Z(n15880));
    LUT4 i2_4_lut_adj_154 (.A(databus[25]), .B(n5_adj_163), .C(n1294[13]), 
         .D(n29544), .Z(n27999)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_154.init = 16'hffec;
    LUT4 select_2068_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1294[4]), 
         .C(rx_data[1]), .D(n29709), .Z(n5_adj_163)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_119)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    PFUMX i9480 (.BLUT(n15885), .ALUT(n28151), .C0(n1747), .Z(n15886));
    LUT4 i2_4_lut_adj_155 (.A(databus[26]), .B(n5_adj_164), .C(n1294[13]), 
         .D(n29545), .Z(n28013)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_155.init = 16'hffec;
    LUT4 select_2068_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1294[4]), 
         .C(rx_data[2]), .D(n29709), .Z(n5_adj_164)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_42_i5_4_lut.init = 16'h88c0;
    PFUMX i13 (.BLUT(n29639), .ALUT(n29766), .C0(n1747), .Z(n29263));
    LUT4 i2_3_lut_rep_299 (.A(n31765), .B(prev_select), .C(n29404), .Z(n31722)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_299.init = 16'h2020;
    LUT4 i1_2_lut_4_lut_adj_156 (.A(n31765), .B(prev_select), .C(n29404), 
         .D(n33447), .Z(n13779)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_156.init = 16'hff20;
    PFUMX i25 (.BLUT(n29808), .ALUT(n29428), .C0(\register_addr[1] ), 
          .Z(n15_adj_123));
    LUT4 i2_4_lut_adj_157 (.A(databus[27]), .B(n5_adj_165), .C(n1294[13]), 
         .D(n29546), .Z(n28023)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_157.init = 16'hffec;
    LUT4 i1_2_lut_rep_417 (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .Z(n31840)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_417.init = 16'heeee;
    LUT4 select_2068_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1294[4]), 
         .C(rx_data[3]), .D(n29709), .Z(n5_adj_165)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_383_3_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(register_addr[5]), .Z(n31806)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_383_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_rep_284_4_lut (.A(n31765), .B(n31826), .C(n29710), .D(prev_select), 
         .Z(n31707)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_rep_284_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_362_3_lut_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(\register_addr[4] ), .D(register_addr[5]), .Z(n31785)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_362_3_lut_4_lut.init = 16'hffef;
    LUT4 i2_4_lut_adj_158 (.A(databus[28]), .B(n5_adj_166), .C(n1294[13]), 
         .D(n29515), .Z(n28026)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_158.init = 16'hffec;
    LUT4 i1_2_lut_rep_384_3_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(\register_addr[3] ), .Z(n31807)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_384_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_159 (.A(n31826), .B(\register_addr[4] ), .C(n29874), 
         .D(n33447), .Z(n14084)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_159.init = 16'hff08;
    LUT4 select_2068_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1294[4]), 
         .C(rx_data[4]), .D(n29709), .Z(n5_adj_166)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_160 (.A(databus[29]), .B(n5_adj_167), .C(n1294[13]), 
         .D(n29520), .Z(n27998)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_160.init = 16'hffec;
    LUT4 i1_2_lut_rep_356_3_lut_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(register_addr[2]), .D(\register_addr[3] ), .Z(n31779)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_356_3_lut_4_lut.init = 16'hfffe;
    LUT4 select_2068_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1294[4]), 
         .C(rx_data[5]), .D(n29709), .Z(n5_adj_167)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_364_3_lut_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(register_addr[5]), .D(\register_addr[3] ), .Z(n31787)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_364_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_371_3_lut_4_lut (.A(register_addr_c[6]), .B(register_addr_c[7]), 
         .C(register_addr[5]), .D(\register_addr[3] ), .Z(n31794)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_371_3_lut_4_lut.init = 16'h0010;
    LUT4 i2_4_lut_adj_161 (.A(databus[30]), .B(n5_adj_168), .C(n1294[13]), 
         .D(n29517), .Z(n28020)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_161.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_adj_162 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [2]), 
         .Z(n29522)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_162.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_163 (.A(\register_addr[4] ), .B(n31763), .C(\read_size[0]_adj_84 ), 
         .Z(n29694)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_163.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_164 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [0]), 
         .Z(n29535)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_164.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_165 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [1]), 
         .Z(n29533)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_165.init = 16'h8080;
    LUT4 reduce_or_455_i1_3_lut (.A(busy), .B(n1294[13]), .C(n1306), .Z(n1405)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_455_i1_3_lut.init = 16'hdcdc;
    LUT4 i1_4_lut_adj_166 (.A(n29627), .B(debug_c_7), .C(n1294[0]), .D(n1294[1]), 
         .Z(n13456)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_166.init = 16'hbbba;
    LUT4 i3_4_lut_adj_167 (.A(sendcount[3]), .B(n31834), .C(sendcount[2]), 
         .D(n31833), .Z(n29627)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_167.init = 16'h0200;
    LUT4 select_2068_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1294[4]), 
         .C(rx_data[6]), .D(n29709), .Z(n5_adj_168)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_168 (.A(databus[31]), .B(n5_adj_170), .C(n1294[13]), 
         .D(n29518), .Z(n28019)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_168.init = 16'hffec;
    LUT4 select_2068_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1294[4]), 
         .C(rx_data[7]), .D(n29709), .Z(n5_adj_170)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2068_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 i15023_3_lut_4_lut (.A(n31757), .B(n1312), .C(n9_adj_74), .D(sendcount[0]), 
         .Z(n18[0])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i15023_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_169 (.A(n31867), .B(n31706), .C(n33447), 
         .D(register_addr[0]), .Z(n13476)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_169.init = 16'hf2f0;
    LUT4 i935_2_lut (.A(n1294[5]), .B(n31783), .Z(n2619)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i935_2_lut.init = 16'h8888;
    LUT4 mux_508_i1_3_lut (.A(n2557), .B(esc_data[0]), .C(n1294[18]), 
         .Z(n2036[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_508_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_170 (.A(n1294[15]), .B(n29860), .C(n30831), .D(n29912), 
         .Z(n2557)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_170.init = 16'h0020;
    LUT4 i23120_2_lut_2_lut (.A(n31783), .B(n9017), .Z(n21320)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i23120_2_lut_2_lut.init = 16'hdddd;
    LUT4 i14790_2_lut (.A(bufcount[0]), .B(n1294[0]), .Z(n15871)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14790_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_adj_171 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [2]), 
         .Z(n29537)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_171.init = 16'h8080;
    LUT4 i1_2_lut_adj_172 (.A(register_addr[0]), .B(\control_reg[7]_adj_85 ), 
         .Z(n8252)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_172.init = 16'h4444;
    LUT4 mux_508_i4_3_lut (.A(n2557), .B(esc_data[3]), .C(n1294[18]), 
         .Z(n2036[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_508_i4_3_lut.init = 16'hcaca;
    LUT4 esc_data_2__bdd_4_lut (.A(esc_data[2]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[4]), .Z(n30831)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam esc_data_2__bdd_4_lut.init = 16'h4801;
    LUT4 i22713_2_lut (.A(esc_data[7]), .B(esc_data[0]), .Z(n29860)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i22713_2_lut.init = 16'hbbbb;
    LUT4 i22765_2_lut (.A(esc_data[5]), .B(esc_data[6]), .Z(n29912)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22765_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_173 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4_adj_86)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_173.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_174 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [3]), 
         .Z(n29538)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_174.init = 16'h8080;
    LUT4 i1_2_lut_adj_175 (.A(register_addr[0]), .B(\control_reg[7]_adj_87 ), 
         .Z(n8261)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_175.init = 16'h4444;
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n31750), .CD(n16067), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_176 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [3]), 
         .Z(n29524)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_176.init = 16'h8080;
    LUT4 i14691_2_lut (.A(sendcount[3]), .B(sendcount[0]), .Z(n17[0])) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i14691_2_lut.init = 16'hdddd;
    LUT4 i2_3_lut_rep_310_4_lut (.A(n31787), .B(n160), .C(\select[4] ), 
         .D(n33446), .Z(n31733)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_310_4_lut.init = 16'h4000;
    LUT4 i14682_2_lut (.A(rx_data[3]), .B(rx_data[1]), .Z(n21052)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14682_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_177 (.A(\register_addr[1] ), .B(\steps_reg[3] ), .Z(n12)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_177.init = 16'h8888;
    LUT4 i15517_3_lut_rep_334 (.A(n1294[13]), .B(n31783), .C(n1312), .Z(n31757)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15517_3_lut_rep_334.init = 16'hc8c8;
    LUT4 i23096_2_lut_rep_305_3_lut (.A(n1294[13]), .B(n31783), .C(n1312), 
         .Z(n31728)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i23096_2_lut_rep_305_3_lut.init = 16'h0808;
    LUT4 i494_2_lut (.A(n1294[3]), .B(n1294[4]), .Z(n1695)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i494_2_lut.init = 16'heeee;
    LUT4 mux_508_i2_3_lut (.A(n2557), .B(esc_data[1]), .C(n1294[18]), 
         .Z(n2036[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_508_i2_3_lut.init = 16'hcaca;
    LUT4 i5463_3_lut (.A(busy), .B(n1306), .C(n1294[19]), .Z(n11867)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5463_3_lut.init = 16'ha8a8;
    LUT4 i23193_4_lut (.A(n7), .B(n29980), .C(n31816), .D(n1294[3]), 
         .Z(n9017)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i23193_4_lut.init = 16'h0544;
    LUT4 i1_2_lut_3_lut_adj_178 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [4]), 
         .Z(n29539)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_178.init = 16'h8080;
    LUT4 mux_1841_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n5613), 
         .Z(n5604[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1841_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_118)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_adj_179 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [5]), 
         .Z(n29540)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_179.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_180 (.A(n31787), .B(\select[4] ), .C(register_addr[2]), 
         .D(\register_addr[4] ), .Z(\arm_select[0] )) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_180.init = 16'h0004;
    LUT4 i1_2_lut_rep_304_4_lut (.A(n31787), .B(\select[4] ), .C(register_addr[2]), 
         .D(\register_addr[4] ), .Z(n31727)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_304_4_lut.init = 16'h0400;
    LUT4 i2_4_lut_adj_181 (.A(n29699), .B(n33446), .C(n31727), .D(prev_select_adj_88), 
         .Z(n3883)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_4_lut_adj_181.init = 16'h0020;
    LUT4 i3_4_lut_adj_182 (.A(n1294[3]), .B(n29473), .C(rx_data[2]), .D(n29623), 
         .Z(n13182)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_182.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_183 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [6]), 
         .Z(n29541)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_183.init = 16'h8080;
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n13568), .CD(n16049), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n13568), .CD(n16049), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n13568), .CD(n16049), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n13568), .CD(n16049), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 i4334_3_lut (.A(n1294[19]), .B(n1294[18]), .C(busy), .Z(n10734)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4334_3_lut.init = 16'hcece;
    LUT4 i1_4_lut_adj_184 (.A(\register_addr[4] ), .B(n2658), .C(n31779), 
         .D(register_addr[5]), .Z(n9089)) /* synthesis lut_function=(A (B)+!A (B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_184.init = 16'hc8cc;
    LUT4 i1_2_lut_3_lut_adj_185 (.A(n1294[3]), .B(n30016), .C(\buffer[4] [7]), 
         .Z(n29542)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_185.init = 16'h8080;
    LUT4 mux_1841_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n5613), 
         .Z(n5604[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1841_i3_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_300_4_lut (.A(\register_addr[4] ), .B(n31794), .C(register_addr[2]), 
         .D(n31826), .Z(n31723)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_300_4_lut.init = 16'h0400;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_116)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_4_lut_adj_186 (.A(\register_addr[4] ), .B(n31794), .C(register_addr[2]), 
         .D(\register_addr[1] ), .Z(n24720)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_186.init = 16'h0004;
    LUT4 mux_1841_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n5613), 
         .Z(n5604[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1841_i2_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_187 (.A(n38), .B(busy), .C(n30674), .D(n1309), 
         .Z(n29123)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_187.init = 16'hfbfa;
    LUT4 i1_2_lut_4_lut_adj_188 (.A(\register_addr[4] ), .B(n31794), .C(register_addr[2]), 
         .D(\register_addr[1] ), .Z(n24690)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_188.init = 16'h0400;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_adj_111)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_adj_189 (.A(n33447), .B(n13606), .Z(n89)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_189.init = 16'heeee;
    LUT4 i1_2_lut_rep_309_4_lut (.A(\register_addr[4] ), .B(n31794), .C(register_addr[2]), 
         .D(\select[4] ), .Z(n31732)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_309_4_lut.init = 16'h0400;
    LUT4 i3_4_lut_adj_190 (.A(n160), .B(prev_select_adj_88), .C(n29404), 
         .D(n31787), .Z(n13606)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i3_4_lut_adj_190.init = 16'h0020;
    LUT4 i22727_4_lut (.A(prev_select_adj_88), .B(register_addr[2]), .C(n29710), 
         .D(n31787), .Z(n29874)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22727_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_191 (.A(n1294[15]), .B(n29860), .C(n30672), .D(n29912), 
         .Z(n38)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_191.init = 16'haaa8;
    LUT4 i1_2_lut_adj_192 (.A(register_addr[0]), .B(rw), .Z(n29710)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_192.init = 16'heeee;
    LUT4 i2_4_lut_adj_193 (.A(n31723), .B(n31773), .C(n33446), .D(prev_select), 
         .Z(n3786)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_193.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_adj_194 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [4]), 
         .Z(n29525)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_194.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_195 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [0]), 
         .Z(n29543)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_195.init = 16'h8080;
    LUT4 i2_3_lut_rep_277_4_lut (.A(\register_addr[1] ), .B(n31779), .C(n185), 
         .D(register_addr[0]), .Z(n31700)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_3_lut_rep_277_4_lut.init = 16'h0010;
    LUT4 i2_3_lut_adj_196 (.A(escape), .B(n4_adj_176), .C(debug_c_7), 
         .Z(n29473)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i2_3_lut_adj_196.init = 16'h4040;
    LUT4 i1_4_lut_adj_197 (.A(rx_data[3]), .B(rx_data[6]), .C(n29632), 
         .D(rx_data[7]), .Z(n4_adj_176)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_197.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_198 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [5]), 
         .Z(n29526)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_198.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_199 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [1]), 
         .Z(n29544)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_199.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_200 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [6]), 
         .Z(n29527)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_200.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_201 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [2]), 
         .Z(n29545)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_201.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_202 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [3]), 
         .Z(n29546)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_202.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_203 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [4]), 
         .Z(n29515)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_203.init = 16'h8080;
    LUT4 i22828_3_lut (.A(n1294[13]), .B(n1294[0]), .C(n1294[4]), .Z(n29980)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22828_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_204 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [5]), 
         .Z(n29520)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_204.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_205 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [6]), 
         .Z(n29517)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_205.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_206 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [7]), 
         .Z(n29528)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_206.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_207 (.A(n1294[3]), .B(n30016), .C(\buffer[5] [7]), 
         .Z(n29518)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_207.init = 16'h8080;
    LUT4 i5462_3_lut (.A(busy), .B(n1309), .C(n1294[16]), .Z(n11865)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5462_3_lut.init = 16'ha8a8;
    LUT4 i14804_2_lut (.A(bufcount[1]), .B(n1294[0]), .Z(n15045)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14804_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_adj_208 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [0]), 
         .Z(n29529)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_208.init = 16'h8080;
    LUT4 i2_3_lut_4_lut_adj_209 (.A(\register_addr[1] ), .B(n31779), .C(n31773), 
         .D(n185), .Z(n3700)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_209.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_210 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [1]), 
         .Z(n29531)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_210.init = 16'h8080;
    LUT4 i2_4_lut_adj_211 (.A(n31779), .B(n185), .C(register_addr[0]), 
         .D(\register_addr[1] ), .Z(n8885)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i2_4_lut_adj_211.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_adj_212 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [2]), 
         .Z(n29521)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_212.init = 16'h8080;
    LUT4 i933_3_lut (.A(n1294[5]), .B(n31783), .C(n1294[10]), .Z(n2617)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i933_3_lut.init = 16'hc8c8;
    LUT4 i1_2_lut_3_lut_adj_213 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [3]), 
         .Z(n29516)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_213.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_214 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [4]), 
         .Z(n29534)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_214.init = 16'h8080;
    LUT4 i5_4_lut (.A(n9_adj_142), .B(n1294[15]), .C(n8_adj_143), .D(n1294[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_215 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [5]), 
         .Z(n29530)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_215.init = 16'h8080;
    LUT4 i1_4_lut_adj_216 (.A(n31823), .B(n1294[18]), .C(n8_adj_177), 
         .D(n1294[6]), .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_216.init = 16'hfffe;
    LUT4 i3_4_lut_adj_217 (.A(n31824), .B(n1294[2]), .C(n4_adj_178), .D(n1294[10]), 
         .Z(n8_adj_177)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_217.init = 16'hfffe;
    LUT4 i1_2_lut_adj_218 (.A(n1294[11]), .B(n1294[7]), .Z(n4_adj_178)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_218.init = 16'heeee;
    LUT4 i4_4_lut (.A(n1294[4]), .B(n29795), .C(n1306), .D(n6_adj_144), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i4_4_lut_adj_219 (.A(n1294[10]), .B(n29795), .C(n31825), .D(n6_adj_179), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_219.init = 16'hfffe;
    LUT4 mux_508_i5_3_lut (.A(n2557), .B(esc_data[4]), .C(n1294[18]), 
         .Z(n2036[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_508_i5_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_220 (.A(n1294[13]), .B(n1294[8]), .Z(n6_adj_179)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_220.init = 16'heeee;
    LUT4 i1_2_lut_rep_294_3_lut_4_lut (.A(\register_addr[4] ), .B(n31787), 
         .C(\register_addr[1] ), .D(register_addr[2]), .Z(n31717)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_294_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_278_4_lut (.A(rw), .B(n31717), .C(prev_select_adj_54), 
         .D(n31827), .Z(n31701)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_278_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_4_lut_adj_221 (.A(\register_addr[4] ), .B(n31787), .C(\register_addr[1] ), 
         .D(register_addr[2]), .Z(n24729)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_221.init = 16'h0100;
    LUT4 i4343_3_lut (.A(n1294[16]), .B(n2557), .C(busy), .Z(n10743)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4343_3_lut.init = 16'hcece;
    LUT4 i1_2_lut_3_lut_adj_222 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [6]), 
         .Z(n29519)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_222.init = 16'h8080;
    LUT4 i1_2_lut_rep_285_3_lut_4_lut (.A(\register_addr[4] ), .B(n31787), 
         .C(n31828), .D(register_addr[2]), .Z(n31708)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_285_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_297_3_lut_4_lut (.A(\register_addr[4] ), .B(n31787), 
         .C(\register_addr[1] ), .D(register_addr[2]), .Z(n31720)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_297_3_lut_4_lut.init = 16'h0010;
    LUT4 n30016_bdd_4_lut_23839 (.A(n30016), .B(n31816), .C(n1294[0]), 
         .D(n1294[3]), .Z(n32223)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n30016_bdd_4_lut_23839.init = 16'hee0f;
    LUT4 i1_2_lut_3_lut_adj_223 (.A(n1294[3]), .B(n30016), .C(\buffer[3] [7]), 
         .Z(n29536)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_223.init = 16'h8080;
    LUT4 i1_2_lut_rep_350 (.A(register_addr[0]), .B(n33447), .Z(n31773)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_350.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_adj_224 (.A(register_addr[0]), .B(n33447), .C(\register_addr[1] ), 
         .Z(n29699)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_224.init = 16'h2020;
    LUT4 i1_2_lut_rep_292_3_lut_4_lut (.A(n160), .B(n31794), .C(prev_select_adj_89), 
         .D(\select[4] ), .Z(n31715)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_292_3_lut_4_lut.init = 16'h0800;
    PFUMX i23766 (.BLUT(n31903), .ALUT(n31904), .C0(sendcount[0]), .Z(n31905));
    LUT4 i1_2_lut_rep_296_3_lut_4_lut (.A(n160), .B(n31794), .C(n33446), 
         .D(\select[4] ), .Z(n31719)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_296_3_lut_4_lut.init = 16'h8000;
    FD1P3AX rw_498_rep_451 (.D(n1294[10]), .SP(n2617), .CK(debug_c_c), 
            .Q(n33446));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_451.GSR = "ENABLED";
    PFUMX i23764 (.BLUT(n31900), .ALUT(n31901), .C0(sendcount[0]), .Z(n31902));
    LUT4 i1_4_lut_adj_225 (.A(n1294[4]), .B(\buffer[0] [0]), .C(n11_adj_99), 
         .D(n14_adj_82), .Z(n28985)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_225.init = 16'heca0;
    PFUMX i23758 (.BLUT(n31891), .ALUT(n31892), .C0(sendcount[0]), .Z(n31893));
    PFUMX i23756 (.BLUT(n31888), .ALUT(n31889), .C0(sendcount[0]), .Z(n31890));
    PFUMX i23754 (.BLUT(n31885), .ALUT(n31886), .C0(n31781), .Z(n31887));
    PFUMX i23752 (.BLUT(n31882), .ALUT(n31883), .C0(sendcount[3]), .Z(n5613));
    PFUMX i23750 (.BLUT(n31879), .ALUT(n31880), .C0(sendcount[0]), .Z(n31881));
    LUT4 i457_2_lut (.A(n5613), .B(n1312), .Z(n1406)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i457_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_226 (.A(n1294[3]), .B(n30016), .C(n1294[13]), 
         .Z(n14_adj_82)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_226.init = 16'hf8f8;
    PFUMX i23748 (.BLUT(n31876), .ALUT(n31877), .C0(sendcount[0]), .Z(n31878));
    LUT4 i1_2_lut_3_lut_adj_227 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [0]), 
         .Z(n29523)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_227.init = 16'h8080;
    PFUMX i23746 (.BLUT(n31873), .ALUT(n31874), .C0(sendcount[0]), .Z(n31875));
    LUT4 i1_2_lut_3_lut_adj_228 (.A(n1294[3]), .B(n30016), .C(\buffer[2] [1]), 
         .Z(n29532)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_228.init = 16'h8080;
    PFUMX i23744 (.BLUT(n31870), .ALUT(n31871), .C0(sendcount[0]), .Z(n31872));
    \UARTTransmitter(baud_div=12)  uart_output (.n33455(n33455), .tx_data({tx_data}), 
            .send(send), .busy(busy), .n31751(n31751), .n31783(n31783), 
            .n10607(n10607), .GND_net(GND_net), .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_c(debug_c_c), .n31783(n31783), 
            .rx_data({rx_data}), .n33455(n33455), .n13070(n13070), .n15(n15), 
            .n10608_c(n10608_c), .debug_c_7(debug_c_7), .n31751(n31751), 
            .n21052(n21052), .n30016(n30016), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (n33455, tx_data, send, busy, 
            n31751, n31783, n10607, GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input n33455;
    input [7:0]tx_data;
    input send;
    output busy;
    input n31751;
    input n31783;
    output n10607;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n30700;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n8997, n2, n30106, n7, n10, n17, n30699, n24391, n31276, 
        n30104, n30105, n31665, n2614, n31664, n14412, n31275, 
        n31752, n29661, n104, n29660, n30698, n4, n29671;
    
    FD1S3IX state__i0 (.D(n30700), .CK(bclk), .CD(n33455), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n8997), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n30106), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15124_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15124_4_lut.init = 16'hfcee;
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 state_1__bdd_4_lut_23525 (.A(state[1]), .B(state[0]), .C(send), 
         .D(state[3]), .Z(n30699)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;
    defparam state_1__bdd_4_lut_23525.init = 16'hb332;
    LUT4 i18071_1_lut (.A(state[3]), .Z(n24391)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i18071_1_lut.init = 16'h5555;
    FD1P3IX busy_34 (.D(n24391), .SP(n31276), .CD(n31751), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 i22951_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n30104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22951_3_lut.init = 16'hcaca;
    LUT4 i22952_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n30105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22952_3_lut.init = 16'hcaca;
    LUT4 send_bdd_4_lut (.A(send), .B(state[3]), .C(state[1]), .D(state[0]), 
         .Z(n31665)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam send_bdd_4_lut.init = 16'h7ffe;
    LUT4 n2613_bdd_4_lut (.A(n31783), .B(state[3]), .C(n2614), .D(state[2]), 
         .Z(n31664)) /* synthesis lut_function=(!((B (D)+!B !(C (D)))+!A)) */ ;
    defparam n2613_bdd_4_lut.init = 16'h2088;
    FD1P3AX state__i3 (.D(n31664), .SP(n14412), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n8997), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n8997), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n8997), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n8997), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n8997), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n8997), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n8997), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 state_2__bdd_4_lut_23799 (.A(send), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n31275)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)))) */ ;
    defparam state_2__bdd_4_lut_23799.init = 16'hc002;
    LUT4 n31275_bdd_2_lut (.A(n31275), .B(state[2]), .Z(n31276)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n31275_bdd_2_lut.init = 16'h2222;
    LUT4 i1_3_lut (.A(state[1]), .B(n31752), .C(state[0]), .Z(n29661)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    LUT4 i1_3_lut_rep_329 (.A(n31783), .B(state[2]), .C(state[3]), .Z(n31752)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut_rep_329.init = 16'h2a2a;
    LUT4 i1_3_lut_4_lut (.A(n31783), .B(state[2]), .C(state[3]), .D(n2614), 
         .Z(n29660)) /* synthesis lut_function=(!((B (C+(D))+!B !(D))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2208;
    PFUMX i23351 (.BLUT(n30699), .ALUT(n30698), .C0(state[2]), .Z(n30700));
    PFUMX i22953 (.BLUT(n30104), .ALUT(n30105), .C0(state[1]), .Z(n30106));
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n31751), .CK(bclk), .Q(n10607)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i2_3_lut_4_lut (.A(n31783), .B(state[2]), .C(n4), .D(n29671), 
         .Z(n8997)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0200;
    FD1P3AX state__i2 (.D(n29660), .SP(n14412), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n29661), .SP(n14412), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 status_led_c_bdd_2_lut_23742_3_lut (.A(n31783), .B(state[2]), .C(n31665), 
         .Z(n14412)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam status_led_c_bdd_2_lut_23742_3_lut.init = 16'hfdfd;
    LUT4 state_1__bdd_2_lut (.A(state[0]), .B(state[3]), .Z(n30698)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 i930_2_lut (.A(state[0]), .B(state[1]), .Z(n2614)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i930_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(send), .B(state[3]), .Z(n29671)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_adj_60 (.A(state[1]), .B(state[0]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_60.init = 16'heeee;
    \ClockDividerP(factor=12)  baud_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .bclk(bclk)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (GND_net, debug_c_c, bclk) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    output bclk;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    
    wire n30210, n49, n56, n50, n16105;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n54, n46, n29866, n52, n42, n48, n34, n27570;
    wire [31:0]n102;
    
    wire n27569, n27568, n27567, n27566, n27565, n27564, n27563, 
        n27562, n27561, n27560, n27559, n27558, n27557, n27556, 
        n27555, n8075, n27618, n27617, n27616, n27615, n27614, 
        n27613, n27612, n27611, n27610, n27609, n27608, n27607, 
        n27606, n27605, n27604, n27603;
    
    LUT4 i23157_4_lut (.A(n30210), .B(n49), .C(n56), .D(n50), .Z(n16105)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23157_4_lut.init = 16'h0002;
    LUT4 i23155_4_lut (.A(count[31]), .B(n54), .C(n46), .D(n29866), 
         .Z(n30210)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23155_4_lut.init = 16'h0100;
    LUT4 i19_4_lut (.A(count[24]), .B(count[27]), .C(count[4]), .D(count[30]), 
         .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(count[5]), .B(n52), .C(n42), .D(count[6]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i20_4_lut (.A(count[7]), .B(count[19]), .C(count[14]), .D(count[22]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(count[16]), .B(n48), .C(n34), .D(count[11]), 
         .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(count[28]), .B(count[2]), .C(count[18]), .D(count[8]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i22719_3_lut (.A(count[3]), .B(count[0]), .C(count[1]), .Z(n29866)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22719_3_lut.init = 16'h8080;
    LUT4 i18_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[21]), .B(count[25]), .Z(n34)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(count[15]), .B(count[29]), .C(count[23]), .D(count[13]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i12_2_lut (.A(count[10]), .B(count[20]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i12_2_lut.init = 16'heeee;
    CCU2D count_2583_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27570), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_33.INIT1 = 16'h0000;
    defparam count_2583_add_4_33.INJECT1_0 = "NO";
    defparam count_2583_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27569), .COUT(n27570), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_31.INJECT1_0 = "NO";
    defparam count_2583_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27568), .COUT(n27569), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_29.INJECT1_0 = "NO";
    defparam count_2583_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27567), .COUT(n27568), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_27.INJECT1_0 = "NO";
    defparam count_2583_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27566), .COUT(n27567), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_25.INJECT1_0 = "NO";
    defparam count_2583_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27565), .COUT(n27566), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_23.INJECT1_0 = "NO";
    defparam count_2583_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27564), .COUT(n27565), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_21.INJECT1_0 = "NO";
    defparam count_2583_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27563), .COUT(n27564), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_19.INJECT1_0 = "NO";
    defparam count_2583_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27562), .COUT(n27563), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_17.INJECT1_0 = "NO";
    defparam count_2583_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27561), .COUT(n27562), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_15.INJECT1_0 = "NO";
    defparam count_2583_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27560), .COUT(n27561), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_13.INJECT1_0 = "NO";
    defparam count_2583_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27559), .COUT(n27560), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_11.INJECT1_0 = "NO";
    defparam count_2583_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27558), .COUT(n27559), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_9.INJECT1_0 = "NO";
    defparam count_2583_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27557), .COUT(n27558), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_7.INJECT1_0 = "NO";
    defparam count_2583_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27556), .COUT(n27557), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_5.INJECT1_0 = "NO";
    defparam count_2583_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27555), .COUT(n27556), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2583_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2583_add_4_3.INJECT1_0 = "NO";
    defparam count_2583_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2583_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27555), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583_add_4_1.INIT0 = 16'hF000;
    defparam count_2583_add_4_1.INIT1 = 16'h0555;
    defparam count_2583_add_4_1.INJECT1_0 = "NO";
    defparam count_2583_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2583__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i0.GSR = "ENABLED";
    FD1S3AX clk_o_14 (.D(n8075), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2583__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i1.GSR = "ENABLED";
    FD1S3IX count_2583__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i2.GSR = "ENABLED";
    FD1S3IX count_2583__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i3.GSR = "ENABLED";
    FD1S3IX count_2583__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i4.GSR = "ENABLED";
    FD1S3IX count_2583__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i5.GSR = "ENABLED";
    FD1S3IX count_2583__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i6.GSR = "ENABLED";
    FD1S3IX count_2583__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i7.GSR = "ENABLED";
    FD1S3IX count_2583__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i8.GSR = "ENABLED";
    FD1S3IX count_2583__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i9.GSR = "ENABLED";
    FD1S3IX count_2583__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i10.GSR = "ENABLED";
    FD1S3IX count_2583__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i11.GSR = "ENABLED";
    FD1S3IX count_2583__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i12.GSR = "ENABLED";
    FD1S3IX count_2583__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i13.GSR = "ENABLED";
    FD1S3IX count_2583__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i14.GSR = "ENABLED";
    FD1S3IX count_2583__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i15.GSR = "ENABLED";
    FD1S3IX count_2583__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i16.GSR = "ENABLED";
    FD1S3IX count_2583__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i17.GSR = "ENABLED";
    FD1S3IX count_2583__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i18.GSR = "ENABLED";
    FD1S3IX count_2583__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i19.GSR = "ENABLED";
    FD1S3IX count_2583__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i20.GSR = "ENABLED";
    FD1S3IX count_2583__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i21.GSR = "ENABLED";
    FD1S3IX count_2583__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i22.GSR = "ENABLED";
    FD1S3IX count_2583__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i23.GSR = "ENABLED";
    FD1S3IX count_2583__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i24.GSR = "ENABLED";
    FD1S3IX count_2583__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i25.GSR = "ENABLED";
    FD1S3IX count_2583__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i26.GSR = "ENABLED";
    FD1S3IX count_2583__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i27.GSR = "ENABLED";
    FD1S3IX count_2583__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i28.GSR = "ENABLED";
    FD1S3IX count_2583__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i29.GSR = "ENABLED";
    FD1S3IX count_2583__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i30.GSR = "ENABLED";
    FD1S3IX count_2583__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16105), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2583__i31.GSR = "ENABLED";
    CCU2D sub_2016_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27618), .S0(n8075));
    defparam sub_2016_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2016_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2016_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2016_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27617), .COUT(n27618));
    defparam sub_2016_add_2_32.INIT0 = 16'h5555;
    defparam sub_2016_add_2_32.INIT1 = 16'h5555;
    defparam sub_2016_add_2_32.INJECT1_0 = "NO";
    defparam sub_2016_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27616), .COUT(n27617));
    defparam sub_2016_add_2_30.INIT0 = 16'h5555;
    defparam sub_2016_add_2_30.INIT1 = 16'h5555;
    defparam sub_2016_add_2_30.INJECT1_0 = "NO";
    defparam sub_2016_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27615), .COUT(n27616));
    defparam sub_2016_add_2_28.INIT0 = 16'h5555;
    defparam sub_2016_add_2_28.INIT1 = 16'h5555;
    defparam sub_2016_add_2_28.INJECT1_0 = "NO";
    defparam sub_2016_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27614), .COUT(n27615));
    defparam sub_2016_add_2_26.INIT0 = 16'h5555;
    defparam sub_2016_add_2_26.INIT1 = 16'h5555;
    defparam sub_2016_add_2_26.INJECT1_0 = "NO";
    defparam sub_2016_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27613), .COUT(n27614));
    defparam sub_2016_add_2_24.INIT0 = 16'h5555;
    defparam sub_2016_add_2_24.INIT1 = 16'h5555;
    defparam sub_2016_add_2_24.INJECT1_0 = "NO";
    defparam sub_2016_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27612), .COUT(n27613));
    defparam sub_2016_add_2_22.INIT0 = 16'h5555;
    defparam sub_2016_add_2_22.INIT1 = 16'h5555;
    defparam sub_2016_add_2_22.INJECT1_0 = "NO";
    defparam sub_2016_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27611), .COUT(n27612));
    defparam sub_2016_add_2_20.INIT0 = 16'h5555;
    defparam sub_2016_add_2_20.INIT1 = 16'h5555;
    defparam sub_2016_add_2_20.INJECT1_0 = "NO";
    defparam sub_2016_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27610), .COUT(n27611));
    defparam sub_2016_add_2_18.INIT0 = 16'h5555;
    defparam sub_2016_add_2_18.INIT1 = 16'h5555;
    defparam sub_2016_add_2_18.INJECT1_0 = "NO";
    defparam sub_2016_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27609), .COUT(n27610));
    defparam sub_2016_add_2_16.INIT0 = 16'h5555;
    defparam sub_2016_add_2_16.INIT1 = 16'h5555;
    defparam sub_2016_add_2_16.INJECT1_0 = "NO";
    defparam sub_2016_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27608), .COUT(n27609));
    defparam sub_2016_add_2_14.INIT0 = 16'h5555;
    defparam sub_2016_add_2_14.INIT1 = 16'h5555;
    defparam sub_2016_add_2_14.INJECT1_0 = "NO";
    defparam sub_2016_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27607), .COUT(n27608));
    defparam sub_2016_add_2_12.INIT0 = 16'h5555;
    defparam sub_2016_add_2_12.INIT1 = 16'h5555;
    defparam sub_2016_add_2_12.INJECT1_0 = "NO";
    defparam sub_2016_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27606), .COUT(n27607));
    defparam sub_2016_add_2_10.INIT0 = 16'h5555;
    defparam sub_2016_add_2_10.INIT1 = 16'h5555;
    defparam sub_2016_add_2_10.INJECT1_0 = "NO";
    defparam sub_2016_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27605), .COUT(n27606));
    defparam sub_2016_add_2_8.INIT0 = 16'h5555;
    defparam sub_2016_add_2_8.INIT1 = 16'h5555;
    defparam sub_2016_add_2_8.INJECT1_0 = "NO";
    defparam sub_2016_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27604), .COUT(n27605));
    defparam sub_2016_add_2_6.INIT0 = 16'h5555;
    defparam sub_2016_add_2_6.INIT1 = 16'h5555;
    defparam sub_2016_add_2_6.INJECT1_0 = "NO";
    defparam sub_2016_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27603), .COUT(n27604));
    defparam sub_2016_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2016_add_2_4.INIT1 = 16'h5555;
    defparam sub_2016_add_2_4.INJECT1_0 = "NO";
    defparam sub_2016_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2016_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27603));
    defparam sub_2016_add_2_2.INIT0 = 16'h0000;
    defparam sub_2016_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2016_add_2_2.INJECT1_0 = "NO";
    defparam sub_2016_add_2_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_c, n31783, rx_data, n33455, 
            n13070, n15, n10608_c, debug_c_7, n31751, n21052, n30016, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31783;
    output [7:0]rx_data;
    input n33455;
    output n13070;
    output n15;
    input n10608_c;
    output debug_c_7;
    input n31751;
    input n21052;
    output n30016;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n8979, n8977, n8975, n8973, n8971, n29005, n8967;
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n272, n192, n212, n8951, n8953, n28753, baud_reset, n30697, 
        n31803, n19, n29780, n13, n13267, n8981, n8983, n8985, 
        n8987, n8989, n8991, n8993, n31821, bclk;
    wire [5:0]n23;
    
    wire n15867, n217, n31836, n10, n31778, n33349, n13255, n28, 
        n13_adj_56, n33347, n33348, n19_adj_57, n31777, n30696, 
        n31801, n29, n15807, n15808, n29075, n15868, n20, n22, 
        n29063;
    wire [7:0]n78;
    
    wire n29071, n33350, n21830, n31837, n4, n21, n30127, n52, 
        n31838, n4_adj_58, n31835, n4_adj_59, n10_adj_60, n26_adj_61, 
        n4_adj_62;
    
    FD1P3AX rdata_i0_i7 (.D(n8979), .SP(n31783), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n8977), .SP(n31783), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n8975), .SP(n31783), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n8973), .SP(n31783), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n8971), .SP(n31783), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n29005), .SP(n31783), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i1 (.D(n8967), .SP(n31783), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(state[3]), .B(rdata[1]), .C(state[2]), .D(n272), 
         .Z(n192)) /* synthesis lut_function=(A (B)+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_4_lut.init = 16'hc8cc;
    LUT4 i1_4_lut_adj_35 (.A(state[2]), .B(rdata[1]), .C(n272), .D(state[3]), 
         .Z(n212)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_4_lut_adj_35.init = 16'hccdc;
    FD1P3AX rdata_i0_i0 (.D(n8951), .SP(n31783), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n8953), .SP(n31783), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n28753), .CK(debug_c_c), .CD(n33455), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n30697), .CK(debug_c_c), .PD(n33455), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n31803), .B(state[0]), .C(state[3]), .D(state[5]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfeff;
    LUT4 i2_4_lut (.A(n29780), .B(rx_data[4]), .C(rx_data[1]), .D(rx_data[3]), 
         .Z(n13070)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'hbfff;
    LUT4 i3_4_lut (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), .D(n29780), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(rx_data[2]), .B(n13), .Z(n29780)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_36 (.A(rdata[1]), .B(rx_data[1]), .C(n13267), .D(n19), 
         .Z(n8981)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_36.init = 16'heca0;
    LUT4 i1_4_lut_adj_37 (.A(rdata[2]), .B(rx_data[2]), .C(n13267), .D(n19), 
         .Z(n8983)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_37.init = 16'heca0;
    LUT4 i1_4_lut_adj_38 (.A(rdata[3]), .B(rx_data[3]), .C(n13267), .D(n19), 
         .Z(n8985)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_38.init = 16'heca0;
    LUT4 i1_4_lut_adj_39 (.A(rdata[4]), .B(rx_data[4]), .C(n13267), .D(n19), 
         .Z(n8987)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_39.init = 16'heca0;
    LUT4 i1_4_lut_adj_40 (.A(rdata[5]), .B(rx_data[5]), .C(n13267), .D(n19), 
         .Z(n8989)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_40.init = 16'heca0;
    LUT4 i1_4_lut_adj_41 (.A(rdata[6]), .B(rx_data[6]), .C(n13267), .D(n19), 
         .Z(n8991)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_41.init = 16'heca0;
    LUT4 i1_4_lut_adj_42 (.A(rdata[7]), .B(rx_data[7]), .C(n13267), .D(n19), 
         .Z(n8993)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_42.init = 16'heca0;
    LUT4 mux_8_i4_3_lut_3_lut (.A(state[3]), .B(n31821), .C(bclk), .Z(n23[3])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam mux_8_i4_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i9461_3_lut_3_lut (.A(state[3]), .B(n31821), .C(bclk), .Z(n15867)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i9461_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i12_3_lut_4_lut (.A(state[5]), .B(n217), .C(state[0]), .D(bclk), 
         .Z(n28753)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i12_3_lut_4_lut.init = 16'hf400;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[4]), .B(n31836), .C(n10608_c), 
         .D(state[3]), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_355_4_lut (.A(state[4]), .B(n31836), .C(state[3]), 
         .D(state[0]), .Z(n31778)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_3_lut_rep_355_4_lut.init = 16'hfffe;
    LUT4 state_0__bdd_2_lut (.A(state[5]), .B(state[4]), .Z(n33349)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam state_0__bdd_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_43 (.A(n13255), .B(rdata[1]), .C(n28), .D(n13_adj_56), 
         .Z(n8967)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_43.init = 16'heca0;
    LUT4 state_4__bdd_3_lut (.A(state[4]), .B(n33347), .C(state[3]), .Z(n33348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam state_4__bdd_3_lut.init = 16'hcaca;
    LUT4 state_3__bdd_4_lut (.A(state[4]), .B(bclk), .C(state[2]), .D(state[1]), 
         .Z(n33347)) /* synthesis lut_function=(A (B+!(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam state_3__bdd_4_lut.init = 16'h9aaa;
    FD1S3IX drdy_51 (.D(n19_adj_57), .CK(debug_c_c), .CD(n31751), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 n10608_c_bdd_4_lut (.A(n10608_c), .B(baud_reset), .C(n31777), 
         .D(state[5]), .Z(n30696)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n10608_c_bdd_4_lut.init = 16'hcfc8;
    LUT4 i3329_3_lut_rep_398 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n31821)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3329_3_lut_rep_398.init = 16'h8080;
    LUT4 i3336_2_lut_rep_378_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n31801)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3336_2_lut_rep_378_4_lut.init = 16'h8000;
    PFUMX i9402 (.BLUT(n29), .ALUT(n15807), .C0(state[0]), .Z(n15808));
    PFUMX i9462 (.BLUT(n29075), .ALUT(n15867), .C0(state[0]), .Z(n15868));
    PFUMX i34 (.BLUT(n20), .ALUT(n22), .C0(state[0]), .Z(n29063));
    LUT4 i1_4_lut_adj_44 (.A(n78[7]), .B(rdata[7]), .C(n13255), .D(n13_adj_56), 
         .Z(n8979)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_44.init = 16'heca0;
    FD1P3AX data_i0_i1 (.D(n8981), .SP(n31783), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n8983), .SP(n31783), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n8985), .SP(n31783), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n8987), .SP(n31783), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n8989), .SP(n31783), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n8991), .SP(n31783), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n8993), .SP(n31783), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n29071), .CK(debug_c_c), .CD(n31751), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n29063), .CK(debug_c_c), .CD(n31751), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n15868), .CK(debug_c_c), .CD(n31751), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n33350), .CK(debug_c_c), .CD(n31751), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n15808), .CK(debug_c_c), .CD(n31751), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    LUT4 i4290_4_lut (.A(rdata[7]), .B(n10608_c), .C(state[2]), .D(n21830), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4290_4_lut.init = 16'hcaaa;
    LUT4 i2_3_lut (.A(state[5]), .B(state[4]), .C(state[0]), .Z(n13255)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i1_4_lut_adj_45 (.A(n78[6]), .B(rdata[6]), .C(n13255), .D(n13_adj_56), 
         .Z(n8977)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_45.init = 16'heca0;
    LUT4 i4292_4_lut (.A(n10608_c), .B(rdata[6]), .C(n31837), .D(n4), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4292_4_lut.init = 16'hccac;
    PFUMX i35 (.BLUT(n21), .ALUT(n30127), .C0(state[0]), .Z(n29071));
    LUT4 i1_2_lut_adj_46 (.A(state[2]), .B(state[1]), .Z(n4)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_adj_46.init = 16'hdddd;
    LUT4 i1_4_lut_adj_47 (.A(n78[5]), .B(rdata[5]), .C(n13255), .D(n13_adj_56), 
         .Z(n8975)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_47.init = 16'heca0;
    LUT4 i4294_4_lut (.A(n10608_c), .B(rdata[5]), .C(state[2]), .D(n21830), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4294_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_48 (.A(n78[4]), .B(rdata[4]), .C(n13255), .D(n13_adj_56), 
         .Z(n8973)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_48.init = 16'heca0;
    LUT4 i4296_4_lut (.A(n10608_c), .B(rdata[4]), .C(n31837), .D(n31836), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4296_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_49 (.A(n13255), .B(rdata[3]), .C(n52), .D(n13_adj_56), 
         .Z(n8971)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_49.init = 16'heca0;
    LUT4 i23170_4_lut (.A(n31838), .B(debug_c_7), .C(n4_adj_58), .D(n31778), 
         .Z(n19_adj_57)) /* synthesis lut_function=(A (B+!(D))+!A (B (C)+!B !((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i23170_4_lut.init = 16'hc8fa;
    LUT4 i18894_4_lut (.A(n31835), .B(n10608_c), .C(rdata[3]), .D(n272), 
         .Z(n52)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B !((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    defparam i18894_4_lut.init = 16'he4f0;
    LUT4 i1_2_lut_rep_412 (.A(state[3]), .B(state[2]), .Z(n31835)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_rep_412.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut (.A(state[3]), .B(state[2]), .C(state[1]), .Z(n4_adj_59)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_rep_413 (.A(state[1]), .B(state[2]), .Z(n31836)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_413.init = 16'heeee;
    PFUMX i18867 (.BLUT(n192), .ALUT(n212), .C0(n10608_c), .Z(n28));
    LUT4 i1_2_lut_rep_354_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .D(state[4]), .Z(n31777)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_354_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_380_3_lut (.A(state[1]), .B(state[2]), .C(state[4]), 
         .Z(n31803)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_380_3_lut.init = 16'hfefe;
    LUT4 i245_2_lut (.A(bclk), .B(state[1]), .Z(n272)) /* synthesis lut_function=(A (B)) */ ;
    defparam i245_2_lut.init = 16'h8888;
    LUT4 i15167_2_lut_rep_414 (.A(bclk), .B(state[3]), .Z(n31837)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15167_2_lut_rep_414.init = 16'h8888;
    LUT4 i1_4_lut_adj_50 (.A(rdata[2]), .B(n13255), .C(n13_adj_56), .D(n10_adj_60), 
         .Z(n29005)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_50.init = 16'heca0;
    LUT4 i15456_2_lut_3_lut (.A(bclk), .B(state[3]), .C(state[1]), .Z(n21830)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15456_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_415 (.A(state[0]), .B(state[5]), .Z(n31838)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_415.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_51 (.A(state[0]), .B(state[5]), .C(state[4]), 
         .Z(n13_adj_56)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_adj_51.init = 16'hefef;
    LUT4 i19_4_lut (.A(n10608_c), .B(rdata[2]), .C(bclk), .D(n4_adj_59), 
         .Z(n10_adj_60)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i19_4_lut.init = 16'hccac;
    LUT4 i22864_4_lut (.A(rx_data[2]), .B(n21052), .C(rx_data[4]), .D(n13), 
         .Z(n30016)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22864_4_lut.init = 16'hfffe;
    PFUMX i24384 (.BLUT(n33349), .ALUT(n33348), .C0(state[0]), .Z(n33350));
    LUT4 i1_4_lut_adj_52 (.A(state[5]), .B(n10), .C(state[1]), .D(n26_adj_61), 
         .Z(n21)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;
    defparam i1_4_lut_adj_52.init = 16'h5111;
    LUT4 i1_3_lut (.A(state[4]), .B(state[2]), .C(state[3]), .Z(n26_adj_61)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i1_3_lut.init = 16'heaea;
    LUT4 i23072_2_lut (.A(state[1]), .B(bclk), .Z(n30127)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i23072_2_lut.init = 16'h9999;
    LUT4 i9401_3_lut_4_lut (.A(state[5]), .B(state[4]), .C(n31801), .D(bclk), 
         .Z(n15807)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(((D)+!C)+!B)) */ ;
    defparam i9401_3_lut_4_lut.init = 16'haa6a;
    LUT4 i3_4_lut_adj_53 (.A(rx_data[5]), .B(rx_data[0]), .C(rx_data[6]), 
         .D(rx_data[7]), .Z(n13)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i3_4_lut_adj_53.init = 16'hfffb;
    LUT4 i1_4_lut_adj_54 (.A(state[5]), .B(n217), .C(n10), .D(n23[3]), 
         .Z(n29075)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_4_lut_adj_54.init = 16'h4505;
    LUT4 n30696_bdd_3_lut (.A(n30696), .B(baud_reset), .C(state[0]), .Z(n30697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30696_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(state[3]), .B(n31803), .C(n10608_c), .D(debug_c_7), 
         .Z(n4_adj_58)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_4_lut_adj_55 (.A(n78[0]), .B(rdata[0]), .C(n13255), .D(n13_adj_56), 
         .Z(n8951)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_55.init = 16'heca0;
    LUT4 i4345_4_lut (.A(n10608_c), .B(rdata[0]), .C(n31836), .D(n4_adj_62), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4345_4_lut.init = 16'hccca;
    LUT4 i1_2_lut_adj_56 (.A(state[3]), .B(bclk), .Z(n4_adj_62)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_adj_56.init = 16'hbbbb;
    LUT4 i2_3_lut_4_lut (.A(state[3]), .B(n31803), .C(state[0]), .D(state[5]), 
         .Z(n13267)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_57 (.A(state[5]), .B(state[2]), .C(n10), .D(n217), 
         .Z(n20)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_57.init = 16'h4505;
    LUT4 i35_3_lut (.A(state[1]), .B(state[2]), .C(bclk), .Z(n22)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i35_3_lut.init = 16'hc6c6;
    LUT4 i1_4_lut_adj_58 (.A(rdata[0]), .B(rx_data[0]), .C(n13267), .D(n19), 
         .Z(n8953)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_58.init = 16'heca0;
    LUT4 i1_4_lut_adj_59 (.A(state[4]), .B(state[2]), .C(state[1]), .D(state[3]), 
         .Z(n217)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_4_lut_adj_59.init = 16'heaaa;
    LUT4 i18937_4_lut (.A(n23[5]), .B(n10), .C(state[5]), .D(n217), 
         .Z(n29)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i18937_4_lut.init = 16'h3a30;
    LUT4 mux_8_i6_3_lut_4_lut (.A(state[5]), .B(state[4]), .C(n31801), 
         .D(bclk), .Z(n23[5])) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam mux_8_i6_3_lut_4_lut.init = 16'h6aaa;
    \ClockDividerP(factor=12)_U0  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .baud_reset(baud_reset), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (bclk, debug_c_c, baud_reset, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input baud_reset;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n8040, n27542;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n27541, n27540, n2766, n27539, n27538, n27537, n27536, 
        n27535, n27534, n27533, n27532, n27531, n27530, n27529, 
        n27528, n27527, n55, n27818, n56, n52, n44, n35, n54, 
        n48, n36, n46, n32, n50, n40, n27650, n27649, n27648, 
        n27647, n27646, n27645, n27644, n27643, n27642, n27641, 
        n27640, n27639, n27638, n27637, n27636, n27635;
    
    FD1S3IX clk_o_14 (.D(n8040), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2582_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27542), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_33.INIT1 = 16'h0000;
    defparam count_2582_add_4_33.INJECT1_0 = "NO";
    defparam count_2582_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27541), .COUT(n27542), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_31.INJECT1_0 = "NO";
    defparam count_2582_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27540), .COUT(n27541), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_29.INJECT1_0 = "NO";
    defparam count_2582_add_4_29.INJECT1_1 = "NO";
    FD1S3IX count_2582__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2766), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i0.GSR = "ENABLED";
    CCU2D count_2582_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27539), .COUT(n27540), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_27.INJECT1_0 = "NO";
    defparam count_2582_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27538), .COUT(n27539), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_25.INJECT1_0 = "NO";
    defparam count_2582_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27537), .COUT(n27538), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_23.INJECT1_0 = "NO";
    defparam count_2582_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27536), .COUT(n27537), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_21.INJECT1_0 = "NO";
    defparam count_2582_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27535), .COUT(n27536), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_19.INJECT1_0 = "NO";
    defparam count_2582_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27534), .COUT(n27535), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_17.INJECT1_0 = "NO";
    defparam count_2582_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27533), .COUT(n27534), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_15.INJECT1_0 = "NO";
    defparam count_2582_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27532), .COUT(n27533), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_13.INJECT1_0 = "NO";
    defparam count_2582_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27531), .COUT(n27532), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_11.INJECT1_0 = "NO";
    defparam count_2582_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27530), .COUT(n27531), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_9.INJECT1_0 = "NO";
    defparam count_2582_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27529), .COUT(n27530), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_7.INJECT1_0 = "NO";
    defparam count_2582_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27528), .COUT(n27529), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_5.INJECT1_0 = "NO";
    defparam count_2582_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27527), .COUT(n27528), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2582_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2582_add_4_3.INJECT1_0 = "NO";
    defparam count_2582_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2582_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27527), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582_add_4_1.INIT0 = 16'hF000;
    defparam count_2582_add_4_1.INIT1 = 16'h0555;
    defparam count_2582_add_4_1.INJECT1_0 = "NO";
    defparam count_2582_add_4_1.INJECT1_1 = "NO";
    LUT4 i1082_4_lut (.A(n55), .B(baud_reset), .C(n27818), .D(n56), 
         .Z(n2766)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i1082_4_lut.init = 16'hccdc;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(count[1]), .B(count[3]), .C(count[0]), .Z(n27818)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    CCU2D sub_2014_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27650), .S0(n8040));
    defparam sub_2014_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2014_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2014_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2014_add_2_cout.INJECT1_1 = "NO";
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i21_4_lut.init = 16'hfffe;
    CCU2D sub_2014_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27649), .COUT(n27650));
    defparam sub_2014_add_2_32.INIT0 = 16'h5555;
    defparam sub_2014_add_2_32.INIT1 = 16'h5555;
    defparam sub_2014_add_2_32.INJECT1_0 = "NO";
    defparam sub_2014_add_2_32.INJECT1_1 = "NO";
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_2_lut.init = 16'heeee;
    CCU2D sub_2014_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27648), .COUT(n27649));
    defparam sub_2014_add_2_30.INIT0 = 16'h5555;
    defparam sub_2014_add_2_30.INIT1 = 16'h5555;
    defparam sub_2014_add_2_30.INJECT1_0 = "NO";
    defparam sub_2014_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27647), .COUT(n27648));
    defparam sub_2014_add_2_28.INIT0 = 16'h5555;
    defparam sub_2014_add_2_28.INIT1 = 16'h5555;
    defparam sub_2014_add_2_28.INJECT1_0 = "NO";
    defparam sub_2014_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27646), .COUT(n27647));
    defparam sub_2014_add_2_26.INIT0 = 16'h5555;
    defparam sub_2014_add_2_26.INIT1 = 16'h5555;
    defparam sub_2014_add_2_26.INJECT1_0 = "NO";
    defparam sub_2014_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27645), .COUT(n27646));
    defparam sub_2014_add_2_24.INIT0 = 16'h5555;
    defparam sub_2014_add_2_24.INIT1 = 16'h5555;
    defparam sub_2014_add_2_24.INJECT1_0 = "NO";
    defparam sub_2014_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27644), .COUT(n27645));
    defparam sub_2014_add_2_22.INIT0 = 16'h5555;
    defparam sub_2014_add_2_22.INIT1 = 16'h5555;
    defparam sub_2014_add_2_22.INJECT1_0 = "NO";
    defparam sub_2014_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27643), .COUT(n27644));
    defparam sub_2014_add_2_20.INIT0 = 16'h5555;
    defparam sub_2014_add_2_20.INIT1 = 16'h5555;
    defparam sub_2014_add_2_20.INJECT1_0 = "NO";
    defparam sub_2014_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27642), .COUT(n27643));
    defparam sub_2014_add_2_18.INIT0 = 16'h5555;
    defparam sub_2014_add_2_18.INIT1 = 16'h5555;
    defparam sub_2014_add_2_18.INJECT1_0 = "NO";
    defparam sub_2014_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27641), .COUT(n27642));
    defparam sub_2014_add_2_16.INIT0 = 16'h5555;
    defparam sub_2014_add_2_16.INIT1 = 16'h5555;
    defparam sub_2014_add_2_16.INJECT1_0 = "NO";
    defparam sub_2014_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27640), .COUT(n27641));
    defparam sub_2014_add_2_14.INIT0 = 16'h5555;
    defparam sub_2014_add_2_14.INIT1 = 16'h5555;
    defparam sub_2014_add_2_14.INJECT1_0 = "NO";
    defparam sub_2014_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27639), .COUT(n27640));
    defparam sub_2014_add_2_12.INIT0 = 16'h5555;
    defparam sub_2014_add_2_12.INIT1 = 16'h5555;
    defparam sub_2014_add_2_12.INJECT1_0 = "NO";
    defparam sub_2014_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27638), .COUT(n27639));
    defparam sub_2014_add_2_10.INIT0 = 16'h5555;
    defparam sub_2014_add_2_10.INIT1 = 16'h5555;
    defparam sub_2014_add_2_10.INJECT1_0 = "NO";
    defparam sub_2014_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27637), .COUT(n27638));
    defparam sub_2014_add_2_8.INIT0 = 16'h5555;
    defparam sub_2014_add_2_8.INIT1 = 16'h5555;
    defparam sub_2014_add_2_8.INJECT1_0 = "NO";
    defparam sub_2014_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27636), .COUT(n27637));
    defparam sub_2014_add_2_6.INIT0 = 16'h5555;
    defparam sub_2014_add_2_6.INIT1 = 16'h5555;
    defparam sub_2014_add_2_6.INJECT1_0 = "NO";
    defparam sub_2014_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27635), .COUT(n27636));
    defparam sub_2014_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2014_add_2_4.INIT1 = 16'h5555;
    defparam sub_2014_add_2_4.INJECT1_0 = "NO";
    defparam sub_2014_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2014_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27635));
    defparam sub_2014_add_2_2.INIT0 = 16'h0000;
    defparam sub_2014_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2014_add_2_2.INJECT1_0 = "NO";
    defparam sub_2014_add_2_2.INJECT1_1 = "NO";
    FD1S3IX count_2582__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2766), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i1.GSR = "ENABLED";
    FD1S3IX count_2582__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2766), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i2.GSR = "ENABLED";
    FD1S3IX count_2582__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2766), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i3.GSR = "ENABLED";
    FD1S3IX count_2582__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2766), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i4.GSR = "ENABLED";
    FD1S3IX count_2582__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2766), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i5.GSR = "ENABLED";
    FD1S3IX count_2582__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2766), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i6.GSR = "ENABLED";
    FD1S3IX count_2582__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2766), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i7.GSR = "ENABLED";
    FD1S3IX count_2582__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2766), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i8.GSR = "ENABLED";
    FD1S3IX count_2582__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2766), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i9.GSR = "ENABLED";
    FD1S3IX count_2582__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i10.GSR = "ENABLED";
    FD1S3IX count_2582__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i11.GSR = "ENABLED";
    FD1S3IX count_2582__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i12.GSR = "ENABLED";
    FD1S3IX count_2582__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i13.GSR = "ENABLED";
    FD1S3IX count_2582__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i14.GSR = "ENABLED";
    FD1S3IX count_2582__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i15.GSR = "ENABLED";
    FD1S3IX count_2582__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i16.GSR = "ENABLED";
    FD1S3IX count_2582__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i17.GSR = "ENABLED";
    FD1S3IX count_2582__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i18.GSR = "ENABLED";
    FD1S3IX count_2582__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i19.GSR = "ENABLED";
    FD1S3IX count_2582__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i20.GSR = "ENABLED";
    FD1S3IX count_2582__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i21.GSR = "ENABLED";
    FD1S3IX count_2582__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i22.GSR = "ENABLED";
    FD1S3IX count_2582__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i23.GSR = "ENABLED";
    FD1S3IX count_2582__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i24.GSR = "ENABLED";
    FD1S3IX count_2582__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i25.GSR = "ENABLED";
    FD1S3IX count_2582__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i26.GSR = "ENABLED";
    FD1S3IX count_2582__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i27.GSR = "ENABLED";
    FD1S3IX count_2582__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i28.GSR = "ENABLED";
    FD1S3IX count_2582__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i29.GSR = "ENABLED";
    FD1S3IX count_2582__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i30.GSR = "ENABLED";
    FD1S3IX count_2582__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2766), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2582__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (read_value, debug_c_c, n2658, 
            VCC_net, GND_net, Stepper_Z_nFault_c, n33450, \read_size[0] , 
            n24720, Stepper_Z_M0_c_0, n13779, n579, prev_step_clk, 
            step_clk, n13757, prev_select, n31732, n31707, n33448, 
            databus, n33449, \control_reg[7] , n31722, Stepper_Z_En_c, 
            Stepper_Z_Dir_c, Stepper_Z_M2_c_2, Stepper_Z_M1_c_1, n27902, 
            n9089, \register_addr[0] , n32, n22, n31711, \register_addr[1] , 
            \read_size[2] , n24690, n33451, n33452, n3786, limit_c_2, 
            n33447, Stepper_Z_Step_c, n8252) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2658;
    input VCC_net;
    input GND_net;
    input Stepper_Z_nFault_c;
    input n33450;
    output \read_size[0] ;
    input n24720;
    output Stepper_Z_M0_c_0;
    input n13779;
    input n579;
    output prev_step_clk;
    output step_clk;
    input n13757;
    output prev_select;
    input n31732;
    input n31707;
    input n33448;
    input [31:0]databus;
    input n33449;
    output \control_reg[7] ;
    input n31722;
    output Stepper_Z_En_c;
    output Stepper_Z_Dir_c;
    output Stepper_Z_M2_c_2;
    output Stepper_Z_M1_c_1;
    output n27902;
    input n9089;
    input \register_addr[0] ;
    input n32;
    input n22;
    input n31711;
    input \register_addr[1] ;
    output \read_size[2] ;
    input n24690;
    input n33451;
    input n33452;
    input n3786;
    input limit_c_2;
    input n33447;
    output Stepper_Z_Step_c;
    input n8252;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n31899, fault_latched;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n3787;
    
    wire limit_latched, n182, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n11634;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n49, n62, n58, n50, n41, n60, n54, n42, n52, n38, 
        n56, n46, n31898, n31897, n27346;
    wire [31:0]n224;
    wire [31:0]n6872;
    
    wire n27345, n27344, n27343, n30055, n30100, n27342, n27341, 
        n27340, n27339, n27338, n27337, n27336, n27335, n27334, 
        n27333, n27332, n27331, n30098, n30099, n29613, n29614, 
        int_step, n30053, n30054;
    wire [7:0]n8251;
    wire [31:0]n6836;
    
    wire n29612;
    
    FD1P3AX read_value__i0 (.D(n31899), .SP(n2658), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3787[0]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n24720), .SP(n2658), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n13779), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13757), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31732), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n31707), .PD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n31707), .PD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n31707), .PD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n31707), .PD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n31707), .CD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n31707), .PD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n31707), .PD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n31707), .PD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n31707), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n31707), .CD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n31707), .CD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n31707), .CD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n31722), .CD(n11634), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n31722), .PD(n33449), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n31722), .PD(n33449), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n31722), .CD(n33449), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n31722), .PD(n33449), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n31722), .CD(n33449), 
            .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n31722), .PD(n33449), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27902)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(steps_reg[9]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(steps_reg[3]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[6]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 n30083_bdd_4_lut_then_4_lut (.A(steps_reg[0]), .B(div_factor_reg[0]), 
         .C(n9089), .D(\register_addr[0] ), .Z(n31898)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam n30083_bdd_4_lut_then_4_lut.init = 16'h0a0c;
    LUT4 n30083_bdd_4_lut_else_4_lut (.A(Stepper_Z_M0_c_0), .B(n9089), .C(limit_latched), 
         .D(\register_addr[0] ), .Z(n31897)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam n30083_bdd_4_lut_else_4_lut.init = 16'h3022;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27346), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    FD1P3IX read_value__i31 (.D(n6872[31]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27345), .COUT(n27346), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27344), .COUT(n27345), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27343), .COUT(n27344), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    FD1P3IX read_value__i28 (.D(n6872[28]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n6872[27]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n6872[26]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n6872[25]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n6872[24]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n6872[23]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n6872[22]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n6872[21]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n6872[20]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n6872[19]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n6872[18]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n6872[17]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n6872[16]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n6872[15]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n6872[14]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n6872[13]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n6872[12]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n6872[11]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n6872[10]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n6872[9]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n6872[8]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6872[7]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6872[6]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6872[5]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6872[4]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6872[3]), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30055), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30100), .SP(n2658), .CD(n9089), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27342), .COUT(n27343), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27341), .COUT(n27342), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27340), .COUT(n27341), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27339), .COUT(n27340), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27338), .COUT(n27339), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27337), .COUT(n27338), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27336), .COUT(n27337), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27335), .COUT(n27336), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27334), .COUT(n27335), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27333), .COUT(n27334), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27332), .COUT(n27333), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27331), .COUT(n27332), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27331), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i22945_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22945_3_lut.init = 16'hcaca;
    LUT4 i22946_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22946_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i29 (.D(n29613), .SP(n2658), .CK(debug_c_c), .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29614), .SP(n2658), .CK(debug_c_c), .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n31711), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i14839_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n6872[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14839_4_lut.init = 16'hc088;
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n13757), .CD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n13757), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n13757), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n13757), .CD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n13757), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n13757), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n13757), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n13757), .CD(n33449), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n13757), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    LUT4 i14840_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n6872[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14840_4_lut.init = 16'hc088;
    LUT4 i14841_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n6872[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14841_4_lut.init = 16'hc088;
    LUT4 i14842_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n6872[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14842_4_lut.init = 16'hc088;
    LUT4 i14843_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n6872[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14843_4_lut.init = 16'hc088;
    FD1P3AX read_size__i2 (.D(n24690), .SP(n2658), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3787[31]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3787[30]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3787[29]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3787[28]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3787[27]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3787[26]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3787[25]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3787[24]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3787[23]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3787[22]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3787[21]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3787[20]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3787[19]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3787[18]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3787[17]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    LUT4 i14844_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n6872[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14844_4_lut.init = 16'hc088;
    FD1S3IX steps_reg__i16 (.D(n3787[16]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3787[15]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3787[14]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3787[13]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3787[12]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3787[11]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3787[10]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3787[9]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3787[8]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3787[7]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3787[6]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3787[5]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3787[4]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3787[3]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3787[2]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3787[1]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i14845_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n6872[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14845_4_lut.init = 16'hc088;
    LUT4 i14846_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n6872[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14846_4_lut.init = 16'hc088;
    LUT4 i14847_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n6872[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14847_4_lut.init = 16'hc088;
    LUT4 i14848_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n6872[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14848_4_lut.init = 16'hc088;
    LUT4 i14849_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n6872[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14849_4_lut.init = 16'hc088;
    LUT4 i14850_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n6872[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14850_4_lut.init = 16'hc088;
    LUT4 i14851_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n6872[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14851_4_lut.init = 16'hc088;
    LUT4 i14852_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n6872[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14852_4_lut.init = 16'hc088;
    LUT4 i14853_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n6872[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14853_4_lut.init = 16'hc088;
    LUT4 i14854_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n6872[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14854_4_lut.init = 16'hc088;
    LUT4 i14855_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n6872[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14855_4_lut.init = 16'hc088;
    LUT4 i14856_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n6872[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14856_4_lut.init = 16'hc088;
    PFUMX i22902 (.BLUT(n30053), .ALUT(n30054), .C0(\register_addr[0] ), 
          .Z(n30055));
    LUT4 i14857_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n6872[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14857_4_lut.init = 16'hc088;
    LUT4 i14858_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n6872[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14858_4_lut.init = 16'hc088;
    LUT4 i14859_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n6872[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14859_4_lut.init = 16'hc088;
    LUT4 i14860_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n6872[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14860_4_lut.init = 16'hc088;
    LUT4 i14838_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8251[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14838_2_lut.init = 16'h2222;
    LUT4 mux_1921_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n6836[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1921_i4_3_lut.init = 16'hcaca;
    LUT4 i14837_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8251[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14837_2_lut.init = 16'h2222;
    LUT4 mux_1921_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n6836[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1921_i5_3_lut.init = 16'hcaca;
    LUT4 i14836_2_lut (.A(Stepper_Z_Dir_c), .B(\register_addr[0] ), .Z(n8251[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14836_2_lut.init = 16'h2222;
    LUT4 mux_1921_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n6836[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1921_i6_3_lut.init = 16'hcaca;
    LUT4 i14835_2_lut (.A(Stepper_Z_En_c), .B(\register_addr[0] ), .Z(n8251[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14835_2_lut.init = 16'h2222;
    LUT4 mux_1921_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n6836[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1921_i7_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(div_factor_reg[29]), .B(n29612), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29613)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(n9089), .Z(n29612)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 mux_1921_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6836[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1921_i8_3_lut.init = 16'hcaca;
    PFUMX i22947 (.BLUT(n30098), .ALUT(n30099), .C0(\register_addr[1] ), 
          .Z(n30100));
    LUT4 i22900_3_lut (.A(Stepper_Z_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22900_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_33 (.A(div_factor_reg[30]), .B(n29612), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29614)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_33.init = 16'hc088;
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    LUT4 i22901_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22901_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n13757), .CD(n33450), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=588, LSE_RLINE=601 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 mux_1521_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3786), 
         .Z(n3787[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3786), 
         .Z(n3787[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3786), 
         .Z(n3787[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3786), 
         .Z(n3787[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3786), 
         .Z(n3787[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3786), 
         .Z(n3787[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3786), 
         .Z(n3787[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3786), 
         .Z(n3787[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3786), 
         .Z(n3787[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3786), 
         .Z(n3787[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3786), 
         .Z(n3787[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3786), 
         .Z(n3787[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3786), 
         .Z(n3787[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3786), 
         .Z(n3787[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3786), 
         .Z(n3787[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3786), 
         .Z(n3787[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3786), 
         .Z(n3787[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3786), 
         .Z(n3787[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3786), 
         .Z(n3787[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3786), 
         .Z(n3787[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3786), 
         .Z(n3787[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3786), 
         .Z(n3787[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3786), .Z(n3787[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3786), .Z(n3787[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3786), .Z(n3787[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3786), .Z(n3787[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3786), .Z(n3787[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3786), .Z(n3787[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3786), .Z(n3787[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3786), .Z(n3787[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3786), .Z(n3787[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1521_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3786), .Z(n3787[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1521_i1_3_lut.init = 16'hcaca;
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    PFUMX mux_1925_i4 (.BLUT(n8251[3]), .ALUT(n6836[3]), .C0(\register_addr[1] ), 
          .Z(n6872[3]));
    PFUMX mux_1925_i5 (.BLUT(n8251[4]), .ALUT(n6836[4]), .C0(\register_addr[1] ), 
          .Z(n6872[4]));
    LUT4 i5234_3_lut (.A(prev_limit_latched), .B(n33447), .C(limit_latched), 
         .Z(n11634)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i5234_3_lut.init = 16'hdcdc;
    PFUMX mux_1925_i6 (.BLUT(n8251[5]), .ALUT(n6836[5]), .C0(\register_addr[1] ), 
          .Z(n6872[5]));
    PFUMX mux_1925_i7 (.BLUT(n8251[6]), .ALUT(n6836[6]), .C0(\register_addr[1] ), 
          .Z(n6872[6]));
    LUT4 i1_2_lut_adj_34 (.A(int_step), .B(control_reg[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_34.init = 16'h9999;
    PFUMX mux_1925_i8 (.BLUT(n8252), .ALUT(n6836[7]), .C0(\register_addr[1] ), 
          .Z(n6872[7]));
    PFUMX i23762 (.BLUT(n31897), .ALUT(n31898), .C0(\register_addr[1] ), 
          .Z(n31899));
    ClockDivider step_clk_gen (.debug_c_c(debug_c_c), .div_factor_reg({div_factor_reg}), 
            .GND_net(GND_net), .step_clk(step_clk), .n33450(n33450), .n33447(n33447)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (debug_c_c, div_factor_reg, GND_net, step_clk, n33450, 
            n33447) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input GND_net;
    output step_clk;
    input n33450;
    input n33447;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n31692, n16111, n27084;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n40;
    
    wire n27085, n27083, n7832, n27082, n7901, n27081, n27080, 
        n27079, n27078, n27077, n27076, n27075, n27074, n27073, 
        n27434;
    wire [31:0]n134;
    
    wire n27433, n27432, n27072, n27431, n27071, n27070, n27069, 
        n27430, n27429, n27068, n27067, n27428, n27427, n27426, 
        n27425, n27424, n27423, n27422, n27421, n27420, n27419, 
        n27114, n7867, n27113, n27112, n27111, n27110, n27109, 
        n27108, n27107, n27106, n27105, n27104, n27103, n27102, 
        n27101, n27100, n27099, n27098, n27097, n27096, n27095, 
        n27094, n27282, n27281, n27093, n27280, n27092, n27091, 
        n27279, n27090, n27089, n27278, n27277, n27276, n27275, 
        n27274, n27273, n27272, n27088, n27271, n27270, n27269, 
        n27268, n27267, n27087, n27086;
    
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2006_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27084), .COUT(n27085));
    defparam sub_2006_add_2_5.INIT0 = 16'h5999;
    defparam sub_2006_add_2_5.INIT1 = 16'h5999;
    defparam sub_2006_add_2_5.INJECT1_0 = "NO";
    defparam sub_2006_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27083), .COUT(n27084));
    defparam sub_2006_add_2_3.INIT0 = 16'h5999;
    defparam sub_2006_add_2_3.INIT1 = 16'h5999;
    defparam sub_2006_add_2_3.INJECT1_0 = "NO";
    defparam sub_2006_add_2_3.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7832), .CK(debug_c_c), .CD(n33450), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2006_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27083));
    defparam sub_2006_add_2_1.INIT0 = 16'h0000;
    defparam sub_2006_add_2_1.INIT1 = 16'h5999;
    defparam sub_2006_add_2_1.INJECT1_0 = "NO";
    defparam sub_2006_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27082), .S1(n7901));
    defparam sub_2007_add_2_33.INIT0 = 16'hf555;
    defparam sub_2007_add_2_33.INIT1 = 16'h0000;
    defparam sub_2007_add_2_33.INJECT1_0 = "NO";
    defparam sub_2007_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27081), .COUT(n27082));
    defparam sub_2007_add_2_31.INIT0 = 16'hf555;
    defparam sub_2007_add_2_31.INIT1 = 16'hf555;
    defparam sub_2007_add_2_31.INJECT1_0 = "NO";
    defparam sub_2007_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27080), .COUT(n27081));
    defparam sub_2007_add_2_29.INIT0 = 16'hf555;
    defparam sub_2007_add_2_29.INIT1 = 16'hf555;
    defparam sub_2007_add_2_29.INJECT1_0 = "NO";
    defparam sub_2007_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27079), .COUT(n27080));
    defparam sub_2007_add_2_27.INIT0 = 16'hf555;
    defparam sub_2007_add_2_27.INIT1 = 16'hf555;
    defparam sub_2007_add_2_27.INJECT1_0 = "NO";
    defparam sub_2007_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27078), .COUT(n27079));
    defparam sub_2007_add_2_25.INIT0 = 16'hf555;
    defparam sub_2007_add_2_25.INIT1 = 16'hf555;
    defparam sub_2007_add_2_25.INJECT1_0 = "NO";
    defparam sub_2007_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27077), .COUT(n27078));
    defparam sub_2007_add_2_23.INIT0 = 16'hf555;
    defparam sub_2007_add_2_23.INIT1 = 16'hf555;
    defparam sub_2007_add_2_23.INJECT1_0 = "NO";
    defparam sub_2007_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27076), .COUT(n27077));
    defparam sub_2007_add_2_21.INIT0 = 16'hf555;
    defparam sub_2007_add_2_21.INIT1 = 16'hf555;
    defparam sub_2007_add_2_21.INJECT1_0 = "NO";
    defparam sub_2007_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27075), .COUT(n27076));
    defparam sub_2007_add_2_19.INIT0 = 16'hf555;
    defparam sub_2007_add_2_19.INIT1 = 16'hf555;
    defparam sub_2007_add_2_19.INJECT1_0 = "NO";
    defparam sub_2007_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27074), .COUT(n27075));
    defparam sub_2007_add_2_17.INIT0 = 16'hf555;
    defparam sub_2007_add_2_17.INIT1 = 16'hf555;
    defparam sub_2007_add_2_17.INJECT1_0 = "NO";
    defparam sub_2007_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27073), .COUT(n27074));
    defparam sub_2007_add_2_15.INIT0 = 16'hf555;
    defparam sub_2007_add_2_15.INIT1 = 16'hf555;
    defparam sub_2007_add_2_15.INJECT1_0 = "NO";
    defparam sub_2007_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27434), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_33.INIT1 = 16'h0000;
    defparam count_2580_add_4_33.INJECT1_0 = "NO";
    defparam count_2580_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27433), .COUT(n27434), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_31.INJECT1_0 = "NO";
    defparam count_2580_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27432), .COUT(n27433), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_29.INJECT1_0 = "NO";
    defparam count_2580_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27072), .COUT(n27073));
    defparam sub_2007_add_2_13.INIT0 = 16'hf555;
    defparam sub_2007_add_2_13.INIT1 = 16'hf555;
    defparam sub_2007_add_2_13.INJECT1_0 = "NO";
    defparam sub_2007_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27431), .COUT(n27432), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_27.INJECT1_0 = "NO";
    defparam count_2580_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27071), .COUT(n27072));
    defparam sub_2007_add_2_11.INIT0 = 16'hf555;
    defparam sub_2007_add_2_11.INIT1 = 16'hf555;
    defparam sub_2007_add_2_11.INJECT1_0 = "NO";
    defparam sub_2007_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27070), .COUT(n27071));
    defparam sub_2007_add_2_9.INIT0 = 16'hf555;
    defparam sub_2007_add_2_9.INIT1 = 16'hf555;
    defparam sub_2007_add_2_9.INJECT1_0 = "NO";
    defparam sub_2007_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27069), .COUT(n27070));
    defparam sub_2007_add_2_7.INIT0 = 16'hf555;
    defparam sub_2007_add_2_7.INIT1 = 16'hf555;
    defparam sub_2007_add_2_7.INJECT1_0 = "NO";
    defparam sub_2007_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27430), .COUT(n27431), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_25.INJECT1_0 = "NO";
    defparam count_2580_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27429), .COUT(n27430), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_23.INJECT1_0 = "NO";
    defparam count_2580_add_4_23.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27068), .COUT(n27069));
    defparam sub_2007_add_2_5.INIT0 = 16'hf555;
    defparam sub_2007_add_2_5.INIT1 = 16'hf555;
    defparam sub_2007_add_2_5.INJECT1_0 = "NO";
    defparam sub_2007_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27067), .COUT(n27068));
    defparam sub_2007_add_2_3.INIT0 = 16'hf555;
    defparam sub_2007_add_2_3.INIT1 = 16'hf555;
    defparam sub_2007_add_2_3.INJECT1_0 = "NO";
    defparam sub_2007_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2007_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27067));
    defparam sub_2007_add_2_1.INIT0 = 16'h0000;
    defparam sub_2007_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2007_add_2_1.INJECT1_0 = "NO";
    defparam sub_2007_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27428), .COUT(n27429), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_21.INJECT1_0 = "NO";
    defparam count_2580_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27427), .COUT(n27428), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_19.INJECT1_0 = "NO";
    defparam count_2580_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27426), .COUT(n27427), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_17.INJECT1_0 = "NO";
    defparam count_2580_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27425), .COUT(n27426), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_15.INJECT1_0 = "NO";
    defparam count_2580_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27424), .COUT(n27425), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_13.INJECT1_0 = "NO";
    defparam count_2580_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27423), .COUT(n27424), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_11.INJECT1_0 = "NO";
    defparam count_2580_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27422), .COUT(n27423), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_9.INJECT1_0 = "NO";
    defparam count_2580_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27421), .COUT(n27422), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_7.INJECT1_0 = "NO";
    defparam count_2580_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27420), .COUT(n27421), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_5.INJECT1_0 = "NO";
    defparam count_2580_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27419), .COUT(n27420), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2580_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2580_add_4_3.INJECT1_0 = "NO";
    defparam count_2580_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2580_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27419), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580_add_4_1.INIT0 = 16'hF000;
    defparam count_2580_add_4_1.INIT1 = 16'h0555;
    defparam count_2580_add_4_1.INJECT1_0 = "NO";
    defparam count_2580_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2580__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i0.GSR = "ENABLED";
    CCU2D sub_2004_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27114), .S1(n7832));
    defparam sub_2004_add_2_33.INIT0 = 16'h5555;
    defparam sub_2004_add_2_33.INIT1 = 16'h0000;
    defparam sub_2004_add_2_33.INJECT1_0 = "NO";
    defparam sub_2004_add_2_33.INJECT1_1 = "NO";
    LUT4 i1009_2_lut_rep_269 (.A(n7867), .B(n33447), .Z(n31692)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1009_2_lut_rep_269.init = 16'heeee;
    CCU2D sub_2004_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27113), .COUT(n27114));
    defparam sub_2004_add_2_31.INIT0 = 16'h5999;
    defparam sub_2004_add_2_31.INIT1 = 16'h5999;
    defparam sub_2004_add_2_31.INJECT1_0 = "NO";
    defparam sub_2004_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27112), .COUT(n27113));
    defparam sub_2004_add_2_29.INIT0 = 16'h5999;
    defparam sub_2004_add_2_29.INIT1 = 16'h5999;
    defparam sub_2004_add_2_29.INJECT1_0 = "NO";
    defparam sub_2004_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27111), .COUT(n27112));
    defparam sub_2004_add_2_27.INIT0 = 16'h5999;
    defparam sub_2004_add_2_27.INIT1 = 16'h5999;
    defparam sub_2004_add_2_27.INJECT1_0 = "NO";
    defparam sub_2004_add_2_27.INJECT1_1 = "NO";
    LUT4 i9705_2_lut_3_lut (.A(n7867), .B(n33447), .C(n7901), .Z(n16111)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9705_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_2004_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27110), .COUT(n27111));
    defparam sub_2004_add_2_25.INIT0 = 16'h5999;
    defparam sub_2004_add_2_25.INIT1 = 16'h5999;
    defparam sub_2004_add_2_25.INJECT1_0 = "NO";
    defparam sub_2004_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27109), .COUT(n27110));
    defparam sub_2004_add_2_23.INIT0 = 16'h5999;
    defparam sub_2004_add_2_23.INIT1 = 16'h5999;
    defparam sub_2004_add_2_23.INJECT1_0 = "NO";
    defparam sub_2004_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27108), .COUT(n27109));
    defparam sub_2004_add_2_21.INIT0 = 16'h5999;
    defparam sub_2004_add_2_21.INIT1 = 16'h5999;
    defparam sub_2004_add_2_21.INJECT1_0 = "NO";
    defparam sub_2004_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27107), .COUT(n27108));
    defparam sub_2004_add_2_19.INIT0 = 16'h5999;
    defparam sub_2004_add_2_19.INIT1 = 16'h5999;
    defparam sub_2004_add_2_19.INJECT1_0 = "NO";
    defparam sub_2004_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27106), .COUT(n27107));
    defparam sub_2004_add_2_17.INIT0 = 16'h5999;
    defparam sub_2004_add_2_17.INIT1 = 16'h5999;
    defparam sub_2004_add_2_17.INJECT1_0 = "NO";
    defparam sub_2004_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27105), .COUT(n27106));
    defparam sub_2004_add_2_15.INIT0 = 16'h5999;
    defparam sub_2004_add_2_15.INIT1 = 16'h5999;
    defparam sub_2004_add_2_15.INJECT1_0 = "NO";
    defparam sub_2004_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27104), .COUT(n27105));
    defparam sub_2004_add_2_13.INIT0 = 16'h5999;
    defparam sub_2004_add_2_13.INIT1 = 16'h5999;
    defparam sub_2004_add_2_13.INJECT1_0 = "NO";
    defparam sub_2004_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27103), .COUT(n27104));
    defparam sub_2004_add_2_11.INIT0 = 16'h5999;
    defparam sub_2004_add_2_11.INIT1 = 16'h5999;
    defparam sub_2004_add_2_11.INJECT1_0 = "NO";
    defparam sub_2004_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27102), .COUT(n27103));
    defparam sub_2004_add_2_9.INIT0 = 16'h5999;
    defparam sub_2004_add_2_9.INIT1 = 16'h5999;
    defparam sub_2004_add_2_9.INJECT1_0 = "NO";
    defparam sub_2004_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27101), .COUT(n27102));
    defparam sub_2004_add_2_7.INIT0 = 16'h5999;
    defparam sub_2004_add_2_7.INIT1 = 16'h5999;
    defparam sub_2004_add_2_7.INJECT1_0 = "NO";
    defparam sub_2004_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27100), .COUT(n27101));
    defparam sub_2004_add_2_5.INIT0 = 16'h5999;
    defparam sub_2004_add_2_5.INIT1 = 16'h5999;
    defparam sub_2004_add_2_5.INJECT1_0 = "NO";
    defparam sub_2004_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27099), .COUT(n27100));
    defparam sub_2004_add_2_3.INIT0 = 16'h5999;
    defparam sub_2004_add_2_3.INIT1 = 16'h5999;
    defparam sub_2004_add_2_3.INJECT1_0 = "NO";
    defparam sub_2004_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2004_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27099));
    defparam sub_2004_add_2_1.INIT0 = 16'h0000;
    defparam sub_2004_add_2_1.INIT1 = 16'h5999;
    defparam sub_2004_add_2_1.INJECT1_0 = "NO";
    defparam sub_2004_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27098), .S1(n7867));
    defparam sub_2006_add_2_33.INIT0 = 16'h5999;
    defparam sub_2006_add_2_33.INIT1 = 16'h0000;
    defparam sub_2006_add_2_33.INJECT1_0 = "NO";
    defparam sub_2006_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27097), .COUT(n27098));
    defparam sub_2006_add_2_31.INIT0 = 16'h5999;
    defparam sub_2006_add_2_31.INIT1 = 16'h5999;
    defparam sub_2006_add_2_31.INJECT1_0 = "NO";
    defparam sub_2006_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    CCU2D sub_2006_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27096), .COUT(n27097));
    defparam sub_2006_add_2_29.INIT0 = 16'h5999;
    defparam sub_2006_add_2_29.INIT1 = 16'h5999;
    defparam sub_2006_add_2_29.INJECT1_0 = "NO";
    defparam sub_2006_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27095), .COUT(n27096));
    defparam sub_2006_add_2_27.INIT0 = 16'h5999;
    defparam sub_2006_add_2_27.INIT1 = 16'h5999;
    defparam sub_2006_add_2_27.INJECT1_0 = "NO";
    defparam sub_2006_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27094), .COUT(n27095));
    defparam sub_2006_add_2_25.INIT0 = 16'h5999;
    defparam sub_2006_add_2_25.INIT1 = 16'h5999;
    defparam sub_2006_add_2_25.INJECT1_0 = "NO";
    defparam sub_2006_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27282), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27281), .COUT(n27282), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27093), .COUT(n27094));
    defparam sub_2006_add_2_23.INIT0 = 16'h5999;
    defparam sub_2006_add_2_23.INIT1 = 16'h5999;
    defparam sub_2006_add_2_23.INJECT1_0 = "NO";
    defparam sub_2006_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27280), .COUT(n27281), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27092), .COUT(n27093));
    defparam sub_2006_add_2_21.INIT0 = 16'h5999;
    defparam sub_2006_add_2_21.INIT1 = 16'h5999;
    defparam sub_2006_add_2_21.INJECT1_0 = "NO";
    defparam sub_2006_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27091), .COUT(n27092));
    defparam sub_2006_add_2_19.INIT0 = 16'h5999;
    defparam sub_2006_add_2_19.INIT1 = 16'h5999;
    defparam sub_2006_add_2_19.INJECT1_0 = "NO";
    defparam sub_2006_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27279), .COUT(n27280), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27090), .COUT(n27091));
    defparam sub_2006_add_2_17.INIT0 = 16'h5999;
    defparam sub_2006_add_2_17.INIT1 = 16'h5999;
    defparam sub_2006_add_2_17.INJECT1_0 = "NO";
    defparam sub_2006_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27089), .COUT(n27090));
    defparam sub_2006_add_2_15.INIT0 = 16'h5999;
    defparam sub_2006_add_2_15.INIT1 = 16'h5999;
    defparam sub_2006_add_2_15.INJECT1_0 = "NO";
    defparam sub_2006_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27278), .COUT(n27279), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27277), .COUT(n27278), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27276), .COUT(n27277), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27275), .COUT(n27276), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27274), .COUT(n27275), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31692), .CD(n16111), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31692), .PD(n16111), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27273), .COUT(n27274), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27272), .COUT(n27273), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    FD1S3IX count_2580__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i1.GSR = "ENABLED";
    FD1S3IX count_2580__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i2.GSR = "ENABLED";
    FD1S3IX count_2580__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i3.GSR = "ENABLED";
    FD1S3IX count_2580__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i4.GSR = "ENABLED";
    FD1S3IX count_2580__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i5.GSR = "ENABLED";
    FD1S3IX count_2580__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i6.GSR = "ENABLED";
    FD1S3IX count_2580__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i7.GSR = "ENABLED";
    FD1S3IX count_2580__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i8.GSR = "ENABLED";
    FD1S3IX count_2580__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i9.GSR = "ENABLED";
    FD1S3IX count_2580__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i10.GSR = "ENABLED";
    FD1S3IX count_2580__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i11.GSR = "ENABLED";
    FD1S3IX count_2580__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i12.GSR = "ENABLED";
    FD1S3IX count_2580__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i13.GSR = "ENABLED";
    FD1S3IX count_2580__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i14.GSR = "ENABLED";
    FD1S3IX count_2580__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i15.GSR = "ENABLED";
    FD1S3IX count_2580__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i16.GSR = "ENABLED";
    FD1S3IX count_2580__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i17.GSR = "ENABLED";
    FD1S3IX count_2580__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i18.GSR = "ENABLED";
    FD1S3IX count_2580__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i19.GSR = "ENABLED";
    FD1S3IX count_2580__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i20.GSR = "ENABLED";
    FD1S3IX count_2580__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i21.GSR = "ENABLED";
    FD1S3IX count_2580__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i22.GSR = "ENABLED";
    FD1S3IX count_2580__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i23.GSR = "ENABLED";
    FD1S3IX count_2580__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i24.GSR = "ENABLED";
    FD1S3IX count_2580__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i25.GSR = "ENABLED";
    FD1S3IX count_2580__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i26.GSR = "ENABLED";
    FD1S3IX count_2580__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i27.GSR = "ENABLED";
    FD1S3IX count_2580__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i28.GSR = "ENABLED";
    FD1S3IX count_2580__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i29.GSR = "ENABLED";
    FD1S3IX count_2580__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i30.GSR = "ENABLED";
    FD1S3IX count_2580__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31692), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2580__i31.GSR = "ENABLED";
    CCU2D sub_2006_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27088), .COUT(n27089));
    defparam sub_2006_add_2_13.INIT0 = 16'h5999;
    defparam sub_2006_add_2_13.INIT1 = 16'h5999;
    defparam sub_2006_add_2_13.INJECT1_0 = "NO";
    defparam sub_2006_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27271), .COUT(n27272), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27270), .COUT(n27271), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27269), .COUT(n27270), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27268), .COUT(n27269), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27267), .COUT(n27268), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27267), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27087), .COUT(n27088));
    defparam sub_2006_add_2_11.INIT0 = 16'h5999;
    defparam sub_2006_add_2_11.INIT1 = 16'h5999;
    defparam sub_2006_add_2_11.INJECT1_0 = "NO";
    defparam sub_2006_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27086), .COUT(n27087));
    defparam sub_2006_add_2_9.INIT0 = 16'h5999;
    defparam sub_2006_add_2_9.INIT1 = 16'h5999;
    defparam sub_2006_add_2_9.INJECT1_0 = "NO";
    defparam sub_2006_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2006_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27085), .COUT(n27086));
    defparam sub_2006_add_2_7.INIT0 = 16'h5999;
    defparam sub_2006_add_2_7.INIT1 = 16'h5999;
    defparam sub_2006_add_2_7.INJECT1_0 = "NO";
    defparam sub_2006_add_2_7.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (\read_size[2] , debug_c_c, n13671, 
            n31720, GND_net, n33451, databus, n3970, n33450, step_clk, 
            n34, prev_step_clk, \read_size[0] , n106, Stepper_X_M0_c_0, 
            n14172, n579, limit_latched, prev_limit_latched, n14124, 
            prev_select, \arm_select[0] , n29552, \register_addr[0] , 
            Stepper_X_M1_c_1, \register_addr[1] , n24, n31713, n31702, 
            n33453, n608, n610, \control_reg[7] , n31701, n10675, 
            Stepper_X_En_c, Stepper_X_Dir_c, Stepper_X_M2_c_2, n27910, 
            VCC_net, Stepper_X_nFault_c, read_value, n31705, limit_c_0, 
            n1, Stepper_X_Step_c, n33447, n33448) /* synthesis syn_module_defined=1 */ ;
    output \read_size[2] ;
    input debug_c_c;
    input n13671;
    input n31720;
    input GND_net;
    input n33451;
    input [31:0]databus;
    input n3970;
    input n33450;
    output step_clk;
    input n34;
    output prev_step_clk;
    output \read_size[0] ;
    input n106;
    output Stepper_X_M0_c_0;
    input n14172;
    input n579;
    output limit_latched;
    output prev_limit_latched;
    input n14124;
    output prev_select;
    input \arm_select[0] ;
    input n29552;
    input \register_addr[0] ;
    output Stepper_X_M1_c_1;
    input \register_addr[1] ;
    input n24;
    input n31713;
    input n31702;
    input n33453;
    input n608;
    input n610;
    output \control_reg[7] ;
    input n31701;
    input n10675;
    output Stepper_X_En_c;
    output Stepper_X_Dir_c;
    output Stepper_X_M2_c_2;
    output n27910;
    input VCC_net;
    input Stepper_X_nFault_c;
    output [31:0]read_value;
    input n31705;
    input limit_c_0;
    input n1;
    output Stepper_X_Step_c;
    input n33447;
    input n33448;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27365;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n224;
    
    wire n27366;
    wire [31:0]n3971;
    
    wire n27364, n27363, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n29554, n29565, fault_latched, n30038, n30039, n30092, 
        n29576, n30093, int_step;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n1_c, n2, n29556, n1_adj_48, n2_adj_49, n29557, n29553, 
        n29558, n1_adj_50, n2_adj_51, n30047, n30048, n30049, n1_adj_52, 
        n2_adj_53, n2_adj_54, n29575, n29574, n29573, n29572, n29571, 
        n29569, n29568, n29567, n29559, n29560, n29570, n29561, 
        n29562, n29563, n29564, n29555, n29566, n49, n62, n58, 
        n50, n30040, n41, n60, n54, n42, n52, n38, n56, n46, 
        n30094;
    wire [31:0]n6278;
    
    wire n27378, n27377, n27376, n27375, n27374, n27373, n27372, 
        n27371, n27370, n27369, n27368, n27367;
    
    FD1P3AX read_size__i2 (.D(n31720), .SP(n13671), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27365), .COUT(n27366), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    FD1S3IX steps_reg__i31 (.D(n3971[31]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    LUT4 mux_1569_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3970), 
         .Z(n3971[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i18_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i30 (.D(n3971[30]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3971[29]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3971[28]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3971[27]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3971[26]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3971[25]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3971[24]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3971[23]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3971[22]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3971[21]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3971[20]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3971[19]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3971[18]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3971[17]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3971[16]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27364), .COUT(n27365), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    FD1S3IX steps_reg__i15 (.D(n3971[15]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3971[14]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3971[13]), .CK(debug_c_c), .CD(n33451), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3971[12]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3971[11]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3971[10]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3971[9]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3971[8]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3971[7]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3971[6]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3971[5]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3971[4]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3971[3]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3971[2]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3971[1]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27363), .COUT(n27364), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n34), .D1(prev_step_clk), 
          .COUT(n27363), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    FD1S3IX steps_reg__i0 (.D(n3971[0]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n106), .SP(n13671), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n14172), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n14124), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    LUT4 mux_1569_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3970), 
         .Z(n3971[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i17_3_lut.init = 16'hcaca;
    FD1S3AX prev_select_174 (.D(\arm_select[0] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(div_factor_reg[21]), .B(n29552), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n29554)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hc088;
    LUT4 mux_1569_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3970), 
         .Z(n3971[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i16_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_10 (.A(div_factor_reg[20]), .B(n29552), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n29565)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_10.init = 16'hc088;
    LUT4 mux_1569_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3970), 
         .Z(n3971[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3970), 
         .Z(n3971[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i14_3_lut.init = 16'hcaca;
    LUT4 i22885_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22885_3_lut.init = 16'hcaca;
    LUT4 i22886_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22886_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3970), 
         .Z(n3971[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3970), 
         .Z(n3971[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3970), 
         .Z(n3971[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3970), 
         .Z(n3971[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i31_3_lut.init = 16'hcaca;
    LUT4 i22939_3_lut (.A(Stepper_X_M0_c_0), .B(div_factor_reg[0]), .C(\register_addr[1] ), 
         .Z(n30092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22939_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_11 (.A(div_factor_reg[19]), .B(n29552), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n29576)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_11.init = 16'hc088;
    LUT4 mux_1569_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3970), 
         .Z(n3971[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i30_3_lut.init = 16'hcaca;
    LUT4 i22940_3_lut (.A(limit_latched), .B(steps_reg[0]), .C(\register_addr[1] ), 
         .Z(n30093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22940_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3970), .Z(n3971[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3970), 
         .Z(n3971[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i29_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n31713), .SP(n24), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i15077_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1_c)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15077_2_lut.init = 16'h2222;
    LUT4 mux_1875_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1875_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_12 (.A(div_factor_reg[18]), .B(n29552), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n29556)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_12.init = 16'hc088;
    LUT4 mux_1569_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3970), 
         .Z(n3971[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3970), .Z(n3971[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i9_3_lut.init = 16'hcaca;
    LUT4 i15076_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_48)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15076_2_lut.init = 16'h2222;
    LUT4 mux_1569_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3970), 
         .Z(n3971[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1875_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2_adj_49)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1875_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_13 (.A(div_factor_reg[17]), .B(n29552), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n29557)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_13.init = 16'hc088;
    LUT4 mux_1569_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3970), .Z(n3971[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_14 (.A(div_factor_reg[16]), .B(n29552), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n29553)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_14.init = 16'hc088;
    LUT4 mux_1569_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3970), .Z(n3971[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3970), 
         .Z(n3971[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3970), .Z(n3971[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i6_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_15 (.A(div_factor_reg[15]), .B(n29552), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n29558)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_15.init = 16'hc088;
    LUT4 mux_1569_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3970), .Z(n3971[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3970), .Z(n3971[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3970), .Z(n3971[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i3_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n31702), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n31702), .PD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n31702), .PD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n31702), .PD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n31702), .PD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n31702), .PD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n31702), .PD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    LUT4 mux_1569_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3970), .Z(n3971[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i2_3_lut.init = 16'hcaca;
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n31702), .PD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n14124), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n14124), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n31701), .CD(n10675), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n31701), .PD(n33453), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n31701), .PD(n33453), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n14172), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n31701), .PD(n33453), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n14172), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n31701), .PD(n33453), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    LUT4 i15071_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_50)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15071_2_lut.init = 16'h2222;
    LUT4 mux_1875_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2_adj_51)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1875_Mux_5_i2_3_lut.init = 16'hcaca;
    PFUMX i22896 (.BLUT(n30047), .ALUT(n30048), .C0(\register_addr[1] ), 
          .Z(n30049));
    LUT4 mux_1569_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3970), 
         .Z(n3971[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i25_3_lut.init = 16'hcaca;
    LUT4 i15070_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_52)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15070_2_lut.init = 16'h2222;
    LUT4 mux_1875_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_53)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1875_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1875_Mux_7_i2_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), 
         .C(\register_addr[0] ), .Z(n2_adj_54)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1875_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1569_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3970), 
         .Z(n3971[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i24_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_16 (.A(div_factor_reg[31]), .B(n29552), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n29575)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_16.init = 16'hc088;
    LUT4 i1_4_lut_adj_17 (.A(div_factor_reg[30]), .B(n29552), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29574)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_17.init = 16'hc088;
    LUT4 i1_4_lut_adj_18 (.A(div_factor_reg[29]), .B(n29552), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29573)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_18.init = 16'hc088;
    LUT4 i1_4_lut_adj_19 (.A(div_factor_reg[28]), .B(n29552), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n29572)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_19.init = 16'hc088;
    LUT4 mux_1569_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3970), 
         .Z(n3971[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i23_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_20 (.A(div_factor_reg[27]), .B(n29552), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n29571)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_20.init = 16'hc088;
    LUT4 i1_4_lut_adj_21 (.A(div_factor_reg[25]), .B(n29552), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n29569)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_21.init = 16'hc088;
    LUT4 i1_4_lut_adj_22 (.A(div_factor_reg[24]), .B(n29552), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n29568)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_22.init = 16'hc088;
    LUT4 i1_4_lut_adj_23 (.A(div_factor_reg[23]), .B(n29552), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n29567)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_23.init = 16'hc088;
    LUT4 i1_4_lut_adj_24 (.A(div_factor_reg[14]), .B(n29552), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n29559)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_24.init = 16'hc088;
    LUT4 i1_4_lut_adj_25 (.A(div_factor_reg[13]), .B(n29552), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n29560)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_25.init = 16'hc088;
    LUT4 i1_4_lut_adj_26 (.A(div_factor_reg[26]), .B(n29552), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n29570)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_26.init = 16'hc088;
    LUT4 i1_4_lut_adj_27 (.A(div_factor_reg[12]), .B(n29552), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n29561)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_27.init = 16'hc088;
    LUT4 i1_4_lut_adj_28 (.A(div_factor_reg[11]), .B(n29552), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n29562)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_28.init = 16'hc088;
    LUT4 mux_1569_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3970), 
         .Z(n3971[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i22_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_29 (.A(div_factor_reg[10]), .B(n29552), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n29563)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_29.init = 16'hc088;
    LUT4 i1_4_lut_adj_30 (.A(div_factor_reg[9]), .B(n29552), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n29564)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_30.init = 16'hc088;
    LUT4 i1_4_lut_adj_31 (.A(div_factor_reg[8]), .B(n29552), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29555)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_31.init = 16'hc088;
    LUT4 mux_1569_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3970), 
         .Z(n3971[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i21_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_32 (.A(div_factor_reg[22]), .B(n29552), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n29566)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_32.init = 16'hc088;
    LUT4 mux_1569_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3970), 
         .Z(n3971[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i20_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27910)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[8]), .B(steps_reg[27]), .C(steps_reg[31]), 
         .D(steps_reg[30]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    PFUMX i22887 (.BLUT(n30038), .ALUT(n30039), .C0(\register_addr[1] ), 
          .Z(n30040));
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[15]), .B(n52), .C(n38), .D(steps_reg[11]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[20]), .B(steps_reg[18]), .C(steps_reg[24]), 
         .D(steps_reg[4]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[9]), .B(steps_reg[12]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 mux_1569_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3970), 
         .Z(n3971[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i19_3_lut.init = 16'hcaca;
    LUT4 i28_4_lut (.A(steps_reg[5]), .B(n56), .C(n46), .D(steps_reg[6]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[7]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[16]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[17]), .B(steps_reg[21]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[19]), .B(steps_reg[3]), .C(steps_reg[22]), 
         .D(steps_reg[13]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[10]), .B(steps_reg[14]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[29]), .B(steps_reg[0]), .C(steps_reg[2]), 
         .D(steps_reg[1]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[28]), .B(steps_reg[23]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    PFUMX i22941 (.BLUT(n30092), .ALUT(n30093), .C0(\register_addr[0] ), 
          .Z(n30094));
    PFUMX mux_1875_Mux_3_i3 (.BLUT(n1_c), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n6278[3]));
    PFUMX mux_1875_Mux_4_i3 (.BLUT(n1_adj_48), .ALUT(n2_adj_49), .C0(\register_addr[1] ), 
          .Z(n6278[4]));
    PFUMX mux_1875_Mux_5_i3 (.BLUT(n1_adj_50), .ALUT(n2_adj_51), .C0(\register_addr[1] ), 
          .Z(n6278[5]));
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    LUT4 mux_1569_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3970), .Z(n3971[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n30094), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    PFUMX mux_1875_Mux_6_i3 (.BLUT(n1_adj_52), .ALUT(n2_adj_53), .C0(\register_addr[1] ), 
          .Z(n6278[6]));
    PFUMX mux_1875_Mux_7_i3 (.BLUT(n1), .ALUT(n2_adj_54), .C0(\register_addr[1] ), 
          .Z(n6278[7]));
    LUT4 i22894_3_lut (.A(Stepper_X_M2_c_2), .B(n34), .C(\register_addr[0] ), 
         .Z(n30047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22894_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i31 (.D(n29575), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29574), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29573), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29572), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29571), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29570), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29569), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29568), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29567), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29566), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29554), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29565), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29576), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29556), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29557), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29553), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29558), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i22895_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22895_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i14 (.D(n29559), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29560), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29561), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29562), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29563), .SP(n13671), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29564), .SP(n13671), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29555), .SP(n13671), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6278[7]), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6278[6]), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6278[5]), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6278[4]), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6278[3]), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30049), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30040), .SP(n13671), .CD(n31705), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27378), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27377), .COUT(n27378), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27376), .COUT(n27377), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27375), .COUT(n27376), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    LUT4 mux_1569_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3970), 
         .Z(n3971[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1569_i32_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27374), .COUT(n27375), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27373), .COUT(n27374), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27372), .COUT(n27373), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27371), .COUT(n27372), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27370), .COUT(n27371), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n14124), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n14124), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27369), .COUT(n27370), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27368), .COUT(n27369), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27367), .COUT(n27368), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n14124), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n14124), .CD(n33453), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=558, LSE_RLINE=571 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27366), .COUT(n27367), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    ClockDivider_U8 step_clk_gen (.div_factor_reg({div_factor_reg}), .GND_net(GND_net), 
            .n33447(n33447), .step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n33448(n33448)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (div_factor_reg, GND_net, n33447, step_clk, debug_c_c, 
            n33448) /* synthesis syn_module_defined=1 */ ;
    input [31:0]div_factor_reg;
    input GND_net;
    input n33447;
    output step_clk;
    input debug_c_c;
    input n33448;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27169, n27170, n27168, n27167, n27166, n7659, n31690, 
        n27165, n7693, n16190, n27164, n27163, n7624, n27314;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n27313;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27312, n27210, n27311, n27310, n27309, n27209, n27208, 
        n27207, n27308, n27206, n27205, n27307, n27306, n27305, 
        n27304, n27204, n27203, n27303, n27202, n27302, n27201, 
        n27301, n27300, n27299, n27200, n27199, n27198, n27197, 
        n27196, n27526, n27195, n27194, n27193, n27192, n27191, 
        n27190, n27525, n27524, n27189, n27188, n27187, n27523, 
        n27186, n27522, n27521, n27520, n27519, n27185, n27518, 
        n27517, n27184, n27183, n27516, n27182, n27515, n27514, 
        n27513, n27512, n27511, n27181, n27180, n27179, n27178, 
        n27177, n27176, n27175, n27174, n27173, n27172, n27171;
    
    CCU2D sub_1997_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27169), .COUT(n27170));
    defparam sub_1997_add_2_15.INIT0 = 16'hf555;
    defparam sub_1997_add_2_15.INIT1 = 16'hf555;
    defparam sub_1997_add_2_15.INJECT1_0 = "NO";
    defparam sub_1997_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27168), .COUT(n27169));
    defparam sub_1997_add_2_13.INIT0 = 16'hf555;
    defparam sub_1997_add_2_13.INIT1 = 16'hf555;
    defparam sub_1997_add_2_13.INJECT1_0 = "NO";
    defparam sub_1997_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27167), .COUT(n27168));
    defparam sub_1997_add_2_11.INIT0 = 16'hf555;
    defparam sub_1997_add_2_11.INIT1 = 16'hf555;
    defparam sub_1997_add_2_11.INJECT1_0 = "NO";
    defparam sub_1997_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27166), .COUT(n27167));
    defparam sub_1997_add_2_9.INIT0 = 16'hf555;
    defparam sub_1997_add_2_9.INIT1 = 16'hf555;
    defparam sub_1997_add_2_9.INJECT1_0 = "NO";
    defparam sub_1997_add_2_9.INJECT1_1 = "NO";
    LUT4 i1001_2_lut_rep_267 (.A(n7659), .B(n33447), .Z(n31690)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1001_2_lut_rep_267.init = 16'heeee;
    CCU2D sub_1997_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27165), .COUT(n27166));
    defparam sub_1997_add_2_7.INIT0 = 16'hf555;
    defparam sub_1997_add_2_7.INIT1 = 16'hf555;
    defparam sub_1997_add_2_7.INJECT1_0 = "NO";
    defparam sub_1997_add_2_7.INJECT1_1 = "NO";
    LUT4 i9813_2_lut_3_lut (.A(n7659), .B(n33447), .C(n7693), .Z(n16190)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9813_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_1997_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27164), .COUT(n27165));
    defparam sub_1997_add_2_5.INIT0 = 16'hf555;
    defparam sub_1997_add_2_5.INIT1 = 16'hf555;
    defparam sub_1997_add_2_5.INJECT1_0 = "NO";
    defparam sub_1997_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27163), .COUT(n27164));
    defparam sub_1997_add_2_3.INIT0 = 16'hf555;
    defparam sub_1997_add_2_3.INIT1 = 16'hf555;
    defparam sub_1997_add_2_3.INJECT1_0 = "NO";
    defparam sub_1997_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27163));
    defparam sub_1997_add_2_1.INIT0 = 16'h0000;
    defparam sub_1997_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1997_add_2_1.INJECT1_0 = "NO";
    defparam sub_1997_add_2_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7624), .CK(debug_c_c), .CD(n33448), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27314), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27313), .COUT(n27314), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    FD1S3IX count_2578__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27312), .COUT(n27313), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27210), .S1(n7624));
    defparam sub_1994_add_2_33.INIT0 = 16'h5555;
    defparam sub_1994_add_2_33.INIT1 = 16'h0000;
    defparam sub_1994_add_2_33.INJECT1_0 = "NO";
    defparam sub_1994_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27311), .COUT(n27312), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27310), .COUT(n27311), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27309), .COUT(n27310), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27209), .COUT(n27210));
    defparam sub_1994_add_2_31.INIT0 = 16'h5999;
    defparam sub_1994_add_2_31.INIT1 = 16'h5999;
    defparam sub_1994_add_2_31.INJECT1_0 = "NO";
    defparam sub_1994_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27208), .COUT(n27209));
    defparam sub_1994_add_2_29.INIT0 = 16'h5999;
    defparam sub_1994_add_2_29.INIT1 = 16'h5999;
    defparam sub_1994_add_2_29.INJECT1_0 = "NO";
    defparam sub_1994_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27207), .COUT(n27208));
    defparam sub_1994_add_2_27.INIT0 = 16'h5999;
    defparam sub_1994_add_2_27.INIT1 = 16'h5999;
    defparam sub_1994_add_2_27.INJECT1_0 = "NO";
    defparam sub_1994_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27308), .COUT(n27309), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27206), .COUT(n27207));
    defparam sub_1994_add_2_25.INIT0 = 16'h5999;
    defparam sub_1994_add_2_25.INIT1 = 16'h5999;
    defparam sub_1994_add_2_25.INJECT1_0 = "NO";
    defparam sub_1994_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27205), .COUT(n27206));
    defparam sub_1994_add_2_23.INIT0 = 16'h5999;
    defparam sub_1994_add_2_23.INIT1 = 16'h5999;
    defparam sub_1994_add_2_23.INJECT1_0 = "NO";
    defparam sub_1994_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27307), .COUT(n27308), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27306), .COUT(n27307), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27305), .COUT(n27306), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27304), .COUT(n27305), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27204), .COUT(n27205));
    defparam sub_1994_add_2_21.INIT0 = 16'h5999;
    defparam sub_1994_add_2_21.INIT1 = 16'h5999;
    defparam sub_1994_add_2_21.INJECT1_0 = "NO";
    defparam sub_1994_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27203), .COUT(n27204));
    defparam sub_1994_add_2_19.INIT0 = 16'h5999;
    defparam sub_1994_add_2_19.INIT1 = 16'h5999;
    defparam sub_1994_add_2_19.INJECT1_0 = "NO";
    defparam sub_1994_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27303), .COUT(n27304), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27202), .COUT(n27203));
    defparam sub_1994_add_2_17.INIT0 = 16'h5999;
    defparam sub_1994_add_2_17.INIT1 = 16'h5999;
    defparam sub_1994_add_2_17.INJECT1_0 = "NO";
    defparam sub_1994_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27302), .COUT(n27303), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27201), .COUT(n27202));
    defparam sub_1994_add_2_15.INIT0 = 16'h5999;
    defparam sub_1994_add_2_15.INIT1 = 16'h5999;
    defparam sub_1994_add_2_15.INJECT1_0 = "NO";
    defparam sub_1994_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27301), .COUT(n27302), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27300), .COUT(n27301), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27299), .COUT(n27300), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27299), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27200), .COUT(n27201));
    defparam sub_1994_add_2_13.INIT0 = 16'h5999;
    defparam sub_1994_add_2_13.INIT1 = 16'h5999;
    defparam sub_1994_add_2_13.INJECT1_0 = "NO";
    defparam sub_1994_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27199), .COUT(n27200));
    defparam sub_1994_add_2_11.INIT0 = 16'h5999;
    defparam sub_1994_add_2_11.INIT1 = 16'h5999;
    defparam sub_1994_add_2_11.INJECT1_0 = "NO";
    defparam sub_1994_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27198), .COUT(n27199));
    defparam sub_1994_add_2_9.INIT0 = 16'h5999;
    defparam sub_1994_add_2_9.INIT1 = 16'h5999;
    defparam sub_1994_add_2_9.INJECT1_0 = "NO";
    defparam sub_1994_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27197), .COUT(n27198));
    defparam sub_1994_add_2_7.INIT0 = 16'h5999;
    defparam sub_1994_add_2_7.INIT1 = 16'h5999;
    defparam sub_1994_add_2_7.INJECT1_0 = "NO";
    defparam sub_1994_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27196), .COUT(n27197));
    defparam sub_1994_add_2_5.INIT0 = 16'h5999;
    defparam sub_1994_add_2_5.INIT1 = 16'h5999;
    defparam sub_1994_add_2_5.INJECT1_0 = "NO";
    defparam sub_1994_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27526), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_33.INIT1 = 16'h0000;
    defparam count_2578_add_4_33.INJECT1_0 = "NO";
    defparam count_2578_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27195), .COUT(n27196));
    defparam sub_1994_add_2_3.INIT0 = 16'h5999;
    defparam sub_1994_add_2_3.INIT1 = 16'h5999;
    defparam sub_1994_add_2_3.INJECT1_0 = "NO";
    defparam sub_1994_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1994_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27195));
    defparam sub_1994_add_2_1.INIT0 = 16'h0000;
    defparam sub_1994_add_2_1.INIT1 = 16'h5999;
    defparam sub_1994_add_2_1.INJECT1_0 = "NO";
    defparam sub_1994_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27194), .S1(n7659));
    defparam sub_1996_add_2_33.INIT0 = 16'h5999;
    defparam sub_1996_add_2_33.INIT1 = 16'h0000;
    defparam sub_1996_add_2_33.INJECT1_0 = "NO";
    defparam sub_1996_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27193), .COUT(n27194));
    defparam sub_1996_add_2_31.INIT0 = 16'h5999;
    defparam sub_1996_add_2_31.INIT1 = 16'h5999;
    defparam sub_1996_add_2_31.INJECT1_0 = "NO";
    defparam sub_1996_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27192), .COUT(n27193));
    defparam sub_1996_add_2_29.INIT0 = 16'h5999;
    defparam sub_1996_add_2_29.INIT1 = 16'h5999;
    defparam sub_1996_add_2_29.INJECT1_0 = "NO";
    defparam sub_1996_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27191), .COUT(n27192));
    defparam sub_1996_add_2_27.INIT0 = 16'h5999;
    defparam sub_1996_add_2_27.INIT1 = 16'h5999;
    defparam sub_1996_add_2_27.INJECT1_0 = "NO";
    defparam sub_1996_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27190), .COUT(n27191));
    defparam sub_1996_add_2_25.INIT0 = 16'h5999;
    defparam sub_1996_add_2_25.INIT1 = 16'h5999;
    defparam sub_1996_add_2_25.INJECT1_0 = "NO";
    defparam sub_1996_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27525), .COUT(n27526), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_31.INJECT1_0 = "NO";
    defparam count_2578_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27524), .COUT(n27525), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_29.INJECT1_0 = "NO";
    defparam count_2578_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27189), .COUT(n27190));
    defparam sub_1996_add_2_23.INIT0 = 16'h5999;
    defparam sub_1996_add_2_23.INIT1 = 16'h5999;
    defparam sub_1996_add_2_23.INJECT1_0 = "NO";
    defparam sub_1996_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27188), .COUT(n27189));
    defparam sub_1996_add_2_21.INIT0 = 16'h5999;
    defparam sub_1996_add_2_21.INIT1 = 16'h5999;
    defparam sub_1996_add_2_21.INJECT1_0 = "NO";
    defparam sub_1996_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27187), .COUT(n27188));
    defparam sub_1996_add_2_19.INIT0 = 16'h5999;
    defparam sub_1996_add_2_19.INIT1 = 16'h5999;
    defparam sub_1996_add_2_19.INJECT1_0 = "NO";
    defparam sub_1996_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27523), .COUT(n27524), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_27.INJECT1_0 = "NO";
    defparam count_2578_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27186), .COUT(n27187));
    defparam sub_1996_add_2_17.INIT0 = 16'h5999;
    defparam sub_1996_add_2_17.INIT1 = 16'h5999;
    defparam sub_1996_add_2_17.INJECT1_0 = "NO";
    defparam sub_1996_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27522), .COUT(n27523), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_25.INJECT1_0 = "NO";
    defparam count_2578_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27521), .COUT(n27522), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_23.INJECT1_0 = "NO";
    defparam count_2578_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27520), .COUT(n27521), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_21.INJECT1_0 = "NO";
    defparam count_2578_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27519), .COUT(n27520), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_19.INJECT1_0 = "NO";
    defparam count_2578_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27185), .COUT(n27186));
    defparam sub_1996_add_2_15.INIT0 = 16'h5999;
    defparam sub_1996_add_2_15.INIT1 = 16'h5999;
    defparam sub_1996_add_2_15.INJECT1_0 = "NO";
    defparam sub_1996_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27518), .COUT(n27519), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_17.INJECT1_0 = "NO";
    defparam count_2578_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27517), .COUT(n27518), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_15.INJECT1_0 = "NO";
    defparam count_2578_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27184), .COUT(n27185));
    defparam sub_1996_add_2_13.INIT0 = 16'h5999;
    defparam sub_1996_add_2_13.INIT1 = 16'h5999;
    defparam sub_1996_add_2_13.INJECT1_0 = "NO";
    defparam sub_1996_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27183), .COUT(n27184));
    defparam sub_1996_add_2_11.INIT0 = 16'h5999;
    defparam sub_1996_add_2_11.INIT1 = 16'h5999;
    defparam sub_1996_add_2_11.INJECT1_0 = "NO";
    defparam sub_1996_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27516), .COUT(n27517), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_13.INJECT1_0 = "NO";
    defparam count_2578_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27182), .COUT(n27183));
    defparam sub_1996_add_2_9.INIT0 = 16'h5999;
    defparam sub_1996_add_2_9.INIT1 = 16'h5999;
    defparam sub_1996_add_2_9.INJECT1_0 = "NO";
    defparam sub_1996_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27515), .COUT(n27516), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_11.INJECT1_0 = "NO";
    defparam count_2578_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27514), .COUT(n27515), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_9.INJECT1_0 = "NO";
    defparam count_2578_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27513), .COUT(n27514), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_7.INJECT1_0 = "NO";
    defparam count_2578_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27512), .COUT(n27513), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_5.INJECT1_0 = "NO";
    defparam count_2578_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27511), .COUT(n27512), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2578_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2578_add_4_3.INJECT1_0 = "NO";
    defparam count_2578_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2578_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27511), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578_add_4_1.INIT0 = 16'hF000;
    defparam count_2578_add_4_1.INIT1 = 16'h0555;
    defparam count_2578_add_4_1.INJECT1_0 = "NO";
    defparam count_2578_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27181), .COUT(n27182));
    defparam sub_1996_add_2_7.INIT0 = 16'h5999;
    defparam sub_1996_add_2_7.INIT1 = 16'h5999;
    defparam sub_1996_add_2_7.INJECT1_0 = "NO";
    defparam sub_1996_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27180), .COUT(n27181));
    defparam sub_1996_add_2_5.INIT0 = 16'h5999;
    defparam sub_1996_add_2_5.INIT1 = 16'h5999;
    defparam sub_1996_add_2_5.INJECT1_0 = "NO";
    defparam sub_1996_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27179), .COUT(n27180));
    defparam sub_1996_add_2_3.INIT0 = 16'h5999;
    defparam sub_1996_add_2_3.INIT1 = 16'h5999;
    defparam sub_1996_add_2_3.INJECT1_0 = "NO";
    defparam sub_1996_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1996_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27179));
    defparam sub_1996_add_2_1.INIT0 = 16'h0000;
    defparam sub_1996_add_2_1.INIT1 = 16'h5999;
    defparam sub_1996_add_2_1.INJECT1_0 = "NO";
    defparam sub_1996_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27178), .S1(n7693));
    defparam sub_1997_add_2_33.INIT0 = 16'hf555;
    defparam sub_1997_add_2_33.INIT1 = 16'h0000;
    defparam sub_1997_add_2_33.INJECT1_0 = "NO";
    defparam sub_1997_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27177), .COUT(n27178));
    defparam sub_1997_add_2_31.INIT0 = 16'hf555;
    defparam sub_1997_add_2_31.INIT1 = 16'hf555;
    defparam sub_1997_add_2_31.INJECT1_0 = "NO";
    defparam sub_1997_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27176), .COUT(n27177));
    defparam sub_1997_add_2_29.INIT0 = 16'hf555;
    defparam sub_1997_add_2_29.INIT1 = 16'hf555;
    defparam sub_1997_add_2_29.INJECT1_0 = "NO";
    defparam sub_1997_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27175), .COUT(n27176));
    defparam sub_1997_add_2_27.INIT0 = 16'hf555;
    defparam sub_1997_add_2_27.INIT1 = 16'hf555;
    defparam sub_1997_add_2_27.INJECT1_0 = "NO";
    defparam sub_1997_add_2_27.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31690), .CD(n16190), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31690), .PD(n16190), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1S3IX count_2578__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i1.GSR = "ENABLED";
    FD1S3IX count_2578__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i2.GSR = "ENABLED";
    FD1S3IX count_2578__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i3.GSR = "ENABLED";
    FD1S3IX count_2578__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i4.GSR = "ENABLED";
    FD1S3IX count_2578__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i5.GSR = "ENABLED";
    FD1S3IX count_2578__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i6.GSR = "ENABLED";
    FD1S3IX count_2578__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i7.GSR = "ENABLED";
    FD1S3IX count_2578__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i8.GSR = "ENABLED";
    FD1S3IX count_2578__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i9.GSR = "ENABLED";
    FD1S3IX count_2578__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i10.GSR = "ENABLED";
    FD1S3IX count_2578__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i11.GSR = "ENABLED";
    FD1S3IX count_2578__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i12.GSR = "ENABLED";
    FD1S3IX count_2578__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i13.GSR = "ENABLED";
    FD1S3IX count_2578__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i14.GSR = "ENABLED";
    FD1S3IX count_2578__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i15.GSR = "ENABLED";
    FD1S3IX count_2578__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i16.GSR = "ENABLED";
    FD1S3IX count_2578__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i17.GSR = "ENABLED";
    FD1S3IX count_2578__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i18.GSR = "ENABLED";
    FD1S3IX count_2578__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i19.GSR = "ENABLED";
    FD1S3IX count_2578__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i20.GSR = "ENABLED";
    FD1S3IX count_2578__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i21.GSR = "ENABLED";
    FD1S3IX count_2578__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i22.GSR = "ENABLED";
    FD1S3IX count_2578__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i23.GSR = "ENABLED";
    FD1S3IX count_2578__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i24.GSR = "ENABLED";
    FD1S3IX count_2578__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i25.GSR = "ENABLED";
    FD1S3IX count_2578__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i26.GSR = "ENABLED";
    FD1S3IX count_2578__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i27.GSR = "ENABLED";
    FD1S3IX count_2578__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i28.GSR = "ENABLED";
    FD1S3IX count_2578__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i29.GSR = "ENABLED";
    FD1S3IX count_2578__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i30.GSR = "ENABLED";
    FD1S3IX count_2578__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31690), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2578__i31.GSR = "ENABLED";
    CCU2D sub_1997_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27174), .COUT(n27175));
    defparam sub_1997_add_2_25.INIT0 = 16'hf555;
    defparam sub_1997_add_2_25.INIT1 = 16'hf555;
    defparam sub_1997_add_2_25.INJECT1_0 = "NO";
    defparam sub_1997_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27173), .COUT(n27174));
    defparam sub_1997_add_2_23.INIT0 = 16'hf555;
    defparam sub_1997_add_2_23.INIT1 = 16'hf555;
    defparam sub_1997_add_2_23.INJECT1_0 = "NO";
    defparam sub_1997_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27172), .COUT(n27173));
    defparam sub_1997_add_2_21.INIT0 = 16'hf555;
    defparam sub_1997_add_2_21.INIT1 = 16'hf555;
    defparam sub_1997_add_2_21.INJECT1_0 = "NO";
    defparam sub_1997_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27171), .COUT(n27172));
    defparam sub_1997_add_2_19.INIT0 = 16'hf555;
    defparam sub_1997_add_2_19.INIT1 = 16'hf555;
    defparam sub_1997_add_2_19.INJECT1_0 = "NO";
    defparam sub_1997_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1997_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27170), .COUT(n27171));
    defparam sub_1997_add_2_17.INIT0 = 16'hf555;
    defparam sub_1997_add_2_17.INIT1 = 16'hf555;
    defparam sub_1997_add_2_17.INJECT1_0 = "NO";
    defparam sub_1997_add_2_17.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (n33447, n7485, n30160, n13719, debug_c_c, 
            n241, n30205, n14176, n30191, n14182, n30189, n14183, 
            n30186, n14186, n29930, n9, n30184, n14187, n30182, 
            n27937, n30195, n27933, n30197, n27924, n30216, n27918, 
            n31694, n30218, n27915, n30152, n27912, GND_net) /* synthesis syn_module_defined=1 */ ;
    input n33447;
    output n7485;
    input n30160;
    output n13719;
    input debug_c_c;
    input n241;
    input n30205;
    output n14176;
    input n30191;
    output n14182;
    input n30189;
    output n14183;
    input n30186;
    output n14186;
    input n29930;
    output n9;
    input n30184;
    output n14187;
    input n30182;
    output n27937;
    input n30195;
    output n27933;
    input n30197;
    output n27924;
    input n30216;
    output n27918;
    output n31694;
    input n30218;
    output n27915;
    input n30152;
    output n27912;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire clk_255kHz, n27418;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n2635, n27417, n27416, n27415, n27414, n27413, n27412, 
        n27411, n27410, n27409, n27408, n27407, n27406, n27405, 
        n27404, n27403, n7520, n27665, n27664, n27663, n27662, 
        n27661, n27660, n27659, n27658, n27657, n27656, n27655, 
        n27654, n27653, n27652, n27651, n27634, n27633, n27632, 
        n27631, n27630, n27629, n27628, n27627, n27626, n27625, 
        n27624, n27623, n27622, n27621, n27620, n27619;
    
    LUT4 i23106_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30160), 
         .Z(n13719)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23106_2_lut_4_lut.init = 16'h1000;
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=518, LSE_RLINE=521 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    LUT4 i23151_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30205), 
         .Z(n14176)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23151_2_lut_4_lut.init = 16'h1000;
    LUT4 i23137_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30191), 
         .Z(n14182)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23137_2_lut_4_lut.init = 16'h1000;
    LUT4 i23135_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30189), 
         .Z(n14183)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23135_2_lut_4_lut.init = 16'h1000;
    LUT4 i23132_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30186), 
         .Z(n14186)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23132_2_lut_4_lut.init = 16'h1000;
    LUT4 i3_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n29930), 
         .Z(n9)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i3_2_lut_4_lut.init = 16'h0010;
    LUT4 i23130_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30184), 
         .Z(n14187)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23130_2_lut_4_lut.init = 16'h1000;
    LUT4 i23128_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30182), 
         .Z(n27937)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23128_2_lut_4_lut.init = 16'h1000;
    LUT4 i23141_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30195), 
         .Z(n27933)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23141_2_lut_4_lut.init = 16'h1000;
    LUT4 i23143_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30197), 
         .Z(n27924)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23143_2_lut_4_lut.init = 16'h1000;
    LUT4 i23162_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30216), 
         .Z(n27918)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23162_2_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_rep_271 (.A(n33447), .B(clk_255kHz), .C(n7485), .Z(n31694)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_3_lut_rep_271.init = 16'h1010;
    LUT4 i23164_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30218), 
         .Z(n27915)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23164_2_lut_4_lut.init = 16'h1000;
    LUT4 i23098_2_lut_4_lut (.A(n33447), .B(clk_255kHz), .C(n7485), .D(n30152), 
         .Z(n27912)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23098_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2575_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27418), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_33.INIT1 = 16'h0000;
    defparam count_2575_add_4_33.INJECT1_0 = "NO";
    defparam count_2575_add_4_33.INJECT1_1 = "NO";
    FD1S3IX count_2575__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2635), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i0.GSR = "ENABLED";
    CCU2D count_2575_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27417), .COUT(n27418), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_31.INJECT1_0 = "NO";
    defparam count_2575_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27416), .COUT(n27417), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_29.INJECT1_0 = "NO";
    defparam count_2575_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27415), .COUT(n27416), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_27.INJECT1_0 = "NO";
    defparam count_2575_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27414), .COUT(n27415), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_25.INJECT1_0 = "NO";
    defparam count_2575_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27413), .COUT(n27414), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_23.INJECT1_0 = "NO";
    defparam count_2575_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27412), .COUT(n27413), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_21.INJECT1_0 = "NO";
    defparam count_2575_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27411), .COUT(n27412), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_19.INJECT1_0 = "NO";
    defparam count_2575_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27410), .COUT(n27411), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_17.INJECT1_0 = "NO";
    defparam count_2575_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27409), .COUT(n27410), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_15.INJECT1_0 = "NO";
    defparam count_2575_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27408), .COUT(n27409), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_13.INJECT1_0 = "NO";
    defparam count_2575_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27407), .COUT(n27408), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_11.INJECT1_0 = "NO";
    defparam count_2575_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27406), .COUT(n27407), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_9.INJECT1_0 = "NO";
    defparam count_2575_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27405), .COUT(n27406), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_7.INJECT1_0 = "NO";
    defparam count_2575_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27404), .COUT(n27405), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_5.INJECT1_0 = "NO";
    defparam count_2575_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27403), .COUT(n27404), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2575_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2575_add_4_3.INJECT1_0 = "NO";
    defparam count_2575_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2575_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27403), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575_add_4_1.INIT0 = 16'hF000;
    defparam count_2575_add_4_1.INIT1 = 16'h0555;
    defparam count_2575_add_4_1.INJECT1_0 = "NO";
    defparam count_2575_add_4_1.INJECT1_1 = "NO";
    LUT4 i951_2_lut (.A(n7520), .B(n33447), .Z(n2635)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i951_2_lut.init = 16'heeee;
    CCU2D add_20536_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27665), 
          .S1(n7485));
    defparam add_20536_32.INIT0 = 16'h5555;
    defparam add_20536_32.INIT1 = 16'h0000;
    defparam add_20536_32.INJECT1_0 = "NO";
    defparam add_20536_32.INJECT1_1 = "NO";
    CCU2D add_20536_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27664), .COUT(n27665));
    defparam add_20536_30.INIT0 = 16'h5555;
    defparam add_20536_30.INIT1 = 16'h5555;
    defparam add_20536_30.INJECT1_0 = "NO";
    defparam add_20536_30.INJECT1_1 = "NO";
    CCU2D add_20536_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27663), .COUT(n27664));
    defparam add_20536_28.INIT0 = 16'h5555;
    defparam add_20536_28.INIT1 = 16'h5555;
    defparam add_20536_28.INJECT1_0 = "NO";
    defparam add_20536_28.INJECT1_1 = "NO";
    CCU2D add_20536_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27662), .COUT(n27663));
    defparam add_20536_26.INIT0 = 16'h5555;
    defparam add_20536_26.INIT1 = 16'h5555;
    defparam add_20536_26.INJECT1_0 = "NO";
    defparam add_20536_26.INJECT1_1 = "NO";
    CCU2D add_20536_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27661), .COUT(n27662));
    defparam add_20536_24.INIT0 = 16'h5555;
    defparam add_20536_24.INIT1 = 16'h5555;
    defparam add_20536_24.INJECT1_0 = "NO";
    defparam add_20536_24.INJECT1_1 = "NO";
    CCU2D add_20536_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27660), .COUT(n27661));
    defparam add_20536_22.INIT0 = 16'h5555;
    defparam add_20536_22.INIT1 = 16'h5555;
    defparam add_20536_22.INJECT1_0 = "NO";
    defparam add_20536_22.INJECT1_1 = "NO";
    CCU2D add_20536_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27659), .COUT(n27660));
    defparam add_20536_20.INIT0 = 16'h5555;
    defparam add_20536_20.INIT1 = 16'h5555;
    defparam add_20536_20.INJECT1_0 = "NO";
    defparam add_20536_20.INJECT1_1 = "NO";
    CCU2D add_20536_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27658), .COUT(n27659));
    defparam add_20536_18.INIT0 = 16'h5555;
    defparam add_20536_18.INIT1 = 16'h5555;
    defparam add_20536_18.INJECT1_0 = "NO";
    defparam add_20536_18.INJECT1_1 = "NO";
    CCU2D add_20536_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27657), .COUT(n27658));
    defparam add_20536_16.INIT0 = 16'h5555;
    defparam add_20536_16.INIT1 = 16'h5555;
    defparam add_20536_16.INJECT1_0 = "NO";
    defparam add_20536_16.INJECT1_1 = "NO";
    CCU2D add_20536_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27656), .COUT(n27657));
    defparam add_20536_14.INIT0 = 16'h5555;
    defparam add_20536_14.INIT1 = 16'h5555;
    defparam add_20536_14.INJECT1_0 = "NO";
    defparam add_20536_14.INJECT1_1 = "NO";
    CCU2D add_20536_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27655), .COUT(n27656));
    defparam add_20536_12.INIT0 = 16'h5555;
    defparam add_20536_12.INIT1 = 16'h5555;
    defparam add_20536_12.INJECT1_0 = "NO";
    defparam add_20536_12.INJECT1_1 = "NO";
    CCU2D add_20536_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27654), .COUT(n27655));
    defparam add_20536_10.INIT0 = 16'h5555;
    defparam add_20536_10.INIT1 = 16'h5555;
    defparam add_20536_10.INJECT1_0 = "NO";
    defparam add_20536_10.INJECT1_1 = "NO";
    CCU2D add_20536_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27653), 
          .COUT(n27654));
    defparam add_20536_8.INIT0 = 16'h5555;
    defparam add_20536_8.INIT1 = 16'h5555;
    defparam add_20536_8.INJECT1_0 = "NO";
    defparam add_20536_8.INJECT1_1 = "NO";
    CCU2D add_20536_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27652), 
          .COUT(n27653));
    defparam add_20536_6.INIT0 = 16'h5555;
    defparam add_20536_6.INIT1 = 16'h5555;
    defparam add_20536_6.INJECT1_0 = "NO";
    defparam add_20536_6.INJECT1_1 = "NO";
    CCU2D add_20536_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27651), 
          .COUT(n27652));
    defparam add_20536_4.INIT0 = 16'h5555;
    defparam add_20536_4.INIT1 = 16'h5aaa;
    defparam add_20536_4.INJECT1_0 = "NO";
    defparam add_20536_4.INJECT1_1 = "NO";
    CCU2D add_20536_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27651));
    defparam add_20536_2.INIT0 = 16'h7000;
    defparam add_20536_2.INIT1 = 16'h5aaa;
    defparam add_20536_2.INJECT1_0 = "NO";
    defparam add_20536_2.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27634), .S0(n7520));
    defparam sub_1989_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1989_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1989_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1989_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27633), .COUT(n27634));
    defparam sub_1989_add_2_32.INIT0 = 16'h5555;
    defparam sub_1989_add_2_32.INIT1 = 16'h5555;
    defparam sub_1989_add_2_32.INJECT1_0 = "NO";
    defparam sub_1989_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27632), .COUT(n27633));
    defparam sub_1989_add_2_30.INIT0 = 16'h5555;
    defparam sub_1989_add_2_30.INIT1 = 16'h5555;
    defparam sub_1989_add_2_30.INJECT1_0 = "NO";
    defparam sub_1989_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27631), .COUT(n27632));
    defparam sub_1989_add_2_28.INIT0 = 16'h5555;
    defparam sub_1989_add_2_28.INIT1 = 16'h5555;
    defparam sub_1989_add_2_28.INJECT1_0 = "NO";
    defparam sub_1989_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27630), .COUT(n27631));
    defparam sub_1989_add_2_26.INIT0 = 16'h5555;
    defparam sub_1989_add_2_26.INIT1 = 16'h5555;
    defparam sub_1989_add_2_26.INJECT1_0 = "NO";
    defparam sub_1989_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27629), .COUT(n27630));
    defparam sub_1989_add_2_24.INIT0 = 16'h5555;
    defparam sub_1989_add_2_24.INIT1 = 16'h5555;
    defparam sub_1989_add_2_24.INJECT1_0 = "NO";
    defparam sub_1989_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27628), .COUT(n27629));
    defparam sub_1989_add_2_22.INIT0 = 16'h5555;
    defparam sub_1989_add_2_22.INIT1 = 16'h5555;
    defparam sub_1989_add_2_22.INJECT1_0 = "NO";
    defparam sub_1989_add_2_22.INJECT1_1 = "NO";
    FD1S3IX count_2575__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2635), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i1.GSR = "ENABLED";
    CCU2D sub_1989_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27627), .COUT(n27628));
    defparam sub_1989_add_2_20.INIT0 = 16'h5555;
    defparam sub_1989_add_2_20.INIT1 = 16'h5555;
    defparam sub_1989_add_2_20.INJECT1_0 = "NO";
    defparam sub_1989_add_2_20.INJECT1_1 = "NO";
    FD1S3IX count_2575__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2635), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i2.GSR = "ENABLED";
    FD1S3IX count_2575__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2635), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i3.GSR = "ENABLED";
    FD1S3IX count_2575__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2635), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i4.GSR = "ENABLED";
    FD1S3IX count_2575__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2635), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i5.GSR = "ENABLED";
    FD1S3IX count_2575__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2635), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i6.GSR = "ENABLED";
    FD1S3IX count_2575__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2635), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i7.GSR = "ENABLED";
    FD1S3IX count_2575__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2635), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i8.GSR = "ENABLED";
    FD1S3IX count_2575__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2635), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i9.GSR = "ENABLED";
    FD1S3IX count_2575__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i10.GSR = "ENABLED";
    FD1S3IX count_2575__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i11.GSR = "ENABLED";
    FD1S3IX count_2575__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i12.GSR = "ENABLED";
    FD1S3IX count_2575__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i13.GSR = "ENABLED";
    FD1S3IX count_2575__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i14.GSR = "ENABLED";
    FD1S3IX count_2575__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i15.GSR = "ENABLED";
    FD1S3IX count_2575__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i16.GSR = "ENABLED";
    FD1S3IX count_2575__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i17.GSR = "ENABLED";
    FD1S3IX count_2575__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i18.GSR = "ENABLED";
    FD1S3IX count_2575__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i19.GSR = "ENABLED";
    FD1S3IX count_2575__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i20.GSR = "ENABLED";
    FD1S3IX count_2575__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i21.GSR = "ENABLED";
    FD1S3IX count_2575__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i22.GSR = "ENABLED";
    FD1S3IX count_2575__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i23.GSR = "ENABLED";
    FD1S3IX count_2575__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i24.GSR = "ENABLED";
    FD1S3IX count_2575__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i25.GSR = "ENABLED";
    FD1S3IX count_2575__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i26.GSR = "ENABLED";
    FD1S3IX count_2575__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i27.GSR = "ENABLED";
    FD1S3IX count_2575__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i28.GSR = "ENABLED";
    FD1S3IX count_2575__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i29.GSR = "ENABLED";
    FD1S3IX count_2575__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i30.GSR = "ENABLED";
    FD1S3IX count_2575__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2635), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2575__i31.GSR = "ENABLED";
    CCU2D sub_1989_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27626), .COUT(n27627));
    defparam sub_1989_add_2_18.INIT0 = 16'h5555;
    defparam sub_1989_add_2_18.INIT1 = 16'h5555;
    defparam sub_1989_add_2_18.INJECT1_0 = "NO";
    defparam sub_1989_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27625), .COUT(n27626));
    defparam sub_1989_add_2_16.INIT0 = 16'h5555;
    defparam sub_1989_add_2_16.INIT1 = 16'h5555;
    defparam sub_1989_add_2_16.INJECT1_0 = "NO";
    defparam sub_1989_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27624), .COUT(n27625));
    defparam sub_1989_add_2_14.INIT0 = 16'h5555;
    defparam sub_1989_add_2_14.INIT1 = 16'h5555;
    defparam sub_1989_add_2_14.INJECT1_0 = "NO";
    defparam sub_1989_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27623), .COUT(n27624));
    defparam sub_1989_add_2_12.INIT0 = 16'h5555;
    defparam sub_1989_add_2_12.INIT1 = 16'h5555;
    defparam sub_1989_add_2_12.INJECT1_0 = "NO";
    defparam sub_1989_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27622), .COUT(n27623));
    defparam sub_1989_add_2_10.INIT0 = 16'h5555;
    defparam sub_1989_add_2_10.INIT1 = 16'h5555;
    defparam sub_1989_add_2_10.INJECT1_0 = "NO";
    defparam sub_1989_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27621), .COUT(n27622));
    defparam sub_1989_add_2_8.INIT0 = 16'h5555;
    defparam sub_1989_add_2_8.INIT1 = 16'h5555;
    defparam sub_1989_add_2_8.INJECT1_0 = "NO";
    defparam sub_1989_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27620), .COUT(n27621));
    defparam sub_1989_add_2_6.INIT0 = 16'h5555;
    defparam sub_1989_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_1989_add_2_6.INJECT1_0 = "NO";
    defparam sub_1989_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27619), .COUT(n27620));
    defparam sub_1989_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1989_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_1989_add_2_4.INJECT1_0 = "NO";
    defparam sub_1989_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_1989_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27619));
    defparam sub_1989_add_2_2.INIT0 = 16'h0000;
    defparam sub_1989_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1989_add_2_2.INJECT1_0 = "NO";
    defparam sub_1989_add_2_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module EncoderPeripheral_U11
//

module EncoderPeripheral_U11 (\read_size[0] , n31762, n24748, read_value, 
            n33457, n31717, encoder_la_c, \register_addr[0] , encoder_lb_c, 
            \read_size[2] , n250, encoder_li_c, n33447, clk_10Hz, 
            n31759, n4144, n47, debug_c_c, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input n31762;
    input n24748;
    output [31:0]read_value;
    input n33457;
    input n31717;
    input encoder_la_c;
    input \register_addr[0] ;
    input encoder_lb_c;
    output \read_size[2] ;
    input n250;
    input encoder_li_c;
    input n33447;
    input clk_10Hz;
    output n31759;
    input n4144;
    output n47;
    input debug_c_c;
    input GND_net;
    input VCC_net;
    
    wire n31762 /* synthesis SET_AS_NETWORK=n31762 */ ;
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(57[14:22])
    wire [31:0]n178;
    
    FD1S3AX read_size_i1 (.D(n24748), .CK(n31762), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_size_i1.GSR = "ENABLED";
    FD1S3IX read_value__i31 (.D(\register[1] [31]), .CK(n31762), .CD(n33457), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1S3IX read_value__i30 (.D(\register[1] [30]), .CK(n31762), .CD(n33457), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1S3IX read_value__i29 (.D(\register[1] [29]), .CK(n31762), .CD(n33457), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1S3IX read_value__i28 (.D(\register[1] [28]), .CK(n31762), .CD(n33457), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1S3IX read_value__i27 (.D(\register[1] [27]), .CK(n31762), .CD(n33457), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1S3IX read_value__i26 (.D(\register[1] [26]), .CK(n31762), .CD(n33457), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1S3IX read_value__i25 (.D(\register[1] [25]), .CK(n31762), .CD(n33457), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1S3IX read_value__i24 (.D(\register[1] [24]), .CK(n31762), .CD(n33457), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1S3IX read_value__i23 (.D(\register[1] [23]), .CK(n31762), .CD(n33457), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1S3IX read_value__i22 (.D(\register[1] [22]), .CK(n31762), .CD(n33457), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1S3IX read_value__i21 (.D(\register[1] [21]), .CK(n31762), .CD(n33457), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1S3IX read_value__i20 (.D(\register[1] [20]), .CK(n31762), .CD(n33457), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1S3IX read_value__i19 (.D(\register[1] [19]), .CK(n31762), .CD(n33457), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1S3IX read_value__i18 (.D(\register[1] [18]), .CK(n31762), .CD(n33457), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1S3IX read_value__i17 (.D(\register[1] [17]), .CK(n31762), .CD(n33457), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1S3IX read_value__i16 (.D(\register[1] [16]), .CK(n31762), .CD(n33457), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1S3IX read_value__i15 (.D(\register[1] [15]), .CK(n31762), .CD(n33457), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1S3IX read_value__i14 (.D(\register[1] [14]), .CK(n31762), .CD(n33457), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1S3IX read_value__i13 (.D(\register[1] [13]), .CK(n31762), .CD(n33457), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1S3IX read_value__i12 (.D(\register[1] [12]), .CK(n31762), .CD(n33457), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1S3IX read_value__i11 (.D(\register[1] [11]), .CK(n31762), .CD(n33457), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1S3IX read_value__i10 (.D(\register[1] [10]), .CK(n31762), .CD(n33457), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1S3IX read_value__i9 (.D(\register[1] [9]), .CK(n31762), .CD(n33457), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1S3IX read_value__i8 (.D(\register[1] [8]), .CK(n31762), .CD(n33457), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1S3IX read_value__i7 (.D(\register[1] [7]), .CK(n31762), .CD(n33457), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(\register[1] [6]), .CK(n31762), .CD(n33457), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(\register[1] [5]), .CK(n31762), .CD(n33457), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(\register[1] [4]), .CK(n31762), .CD(n33457), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n178[2]), .CK(n31762), .CD(n31717), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i1 (.D(n178[1]), .CK(n31762), .CD(n31717), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n178[3]), .CK(n31762), .CD(n31717), .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i3.GSR = "ENABLED";
    LUT4 mux_113_Mux_3_i1_3_lut (.A(encoder_la_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n178[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(76[29:42])
    defparam mux_113_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_113_Mux_2_i1_3_lut (.A(encoder_lb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n178[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(76[29:42])
    defparam mux_113_Mux_2_i1_3_lut.init = 16'hcaca;
    FD1S3AX read_size_i2 (.D(n250), .CK(n31762), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_size_i2.GSR = "ENABLED";
    LUT4 mux_113_Mux_1_i1_3_lut (.A(encoder_li_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n178[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(76[29:42])
    defparam mux_113_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 i4_2_lut_rep_336 (.A(n33447), .B(clk_10Hz), .Z(n31759)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(63[18:34])
    defparam i4_2_lut_rep_336.init = 16'heeee;
    LUT4 i15205_2_lut_3_lut (.A(n33447), .B(clk_10Hz), .C(n4144), .Z(n47)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(63[18:34])
    defparam i15205_2_lut_3_lut.init = 16'h1010;
    FD1S3IX read_value__i0 (.D(\register[1] [0]), .CK(n31762), .CD(n33457), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=646, LSE_RLINE=656 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i0.GSR = "ENABLED";
    QuadratureDecoder_U6 q (.\register[1] ({\register[1] }), .debug_c_c(debug_c_c), 
            .n31759(n31759), .encoder_la_c(encoder_la_c), .GND_net(GND_net), 
            .VCC_net(VCC_net), .encoder_lb_c(encoder_lb_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(88[20] 92[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder_U6
//

module QuadratureDecoder_U6 (\register[1] , debug_c_c, n31759, encoder_la_c, 
            GND_net, VCC_net, encoder_lb_c) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[1] ;
    input debug_c_c;
    input n31759;
    input encoder_la_c;
    input GND_net;
    input VCC_net;
    input encoder_lb_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n13565;
    wire [31:0]n100;
    
    wire n27010, quadB_delayed, n27011, n27009, n27008, n27007, 
        n27006, n27005, n27004, n27003, n27002, quadA_delayed, n27017, 
        n27016, n27015, n6, n27014, n27013, n27012;
    
    FD1P3IX count__i0 (.D(n100[0]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX count__i31 (.D(n100[31]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n100[30]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n100[29]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n100[28]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n100[27]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n100[26]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n100[25]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n100[24]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n100[23]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n100[22]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n100[21]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n100[20]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n100[19]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n100[18]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n100[17]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n100[16]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n100[15]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n100[14]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n100[13]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n100[12]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n100[11]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n100[10]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n100[9]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n100[8]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n100[7]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n100[6]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n100[5]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n100[4]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n100[3]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n100[2]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n100[1]), .SP(n13565), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i1.GSR = "ENABLED";
    CCU2D add_1663_19 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [16]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [17]), 
          .D1(GND_net), .CIN(n27010), .COUT(n27011), .S0(n100[16]), 
          .S1(n100[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_19.INIT0 = 16'h6969;
    defparam add_1663_19.INIT1 = 16'h6969;
    defparam add_1663_19.INJECT1_0 = "NO";
    defparam add_1663_19.INJECT1_1 = "NO";
    CCU2D add_1663_17 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [14]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [15]), 
          .D1(GND_net), .CIN(n27009), .COUT(n27010), .S0(n100[14]), 
          .S1(n100[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_17.INIT0 = 16'h6969;
    defparam add_1663_17.INIT1 = 16'h6969;
    defparam add_1663_17.INJECT1_0 = "NO";
    defparam add_1663_17.INJECT1_1 = "NO";
    CCU2D add_1663_15 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [12]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [13]), 
          .D1(GND_net), .CIN(n27008), .COUT(n27009), .S0(n100[12]), 
          .S1(n100[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_15.INIT0 = 16'h6969;
    defparam add_1663_15.INIT1 = 16'h6969;
    defparam add_1663_15.INJECT1_0 = "NO";
    defparam add_1663_15.INJECT1_1 = "NO";
    CCU2D add_1663_13 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [10]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [11]), 
          .D1(GND_net), .CIN(n27007), .COUT(n27008), .S0(n100[10]), 
          .S1(n100[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_13.INIT0 = 16'h6969;
    defparam add_1663_13.INIT1 = 16'h6969;
    defparam add_1663_13.INJECT1_0 = "NO";
    defparam add_1663_13.INJECT1_1 = "NO";
    CCU2D add_1663_11 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [8]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [9]), 
          .D1(GND_net), .CIN(n27006), .COUT(n27007), .S0(n100[8]), .S1(n100[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_11.INIT0 = 16'h6969;
    defparam add_1663_11.INIT1 = 16'h6969;
    defparam add_1663_11.INJECT1_0 = "NO";
    defparam add_1663_11.INJECT1_1 = "NO";
    CCU2D add_1663_9 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [6]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [7]), 
          .D1(GND_net), .CIN(n27005), .COUT(n27006), .S0(n100[6]), .S1(n100[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_9.INIT0 = 16'h6969;
    defparam add_1663_9.INIT1 = 16'h6969;
    defparam add_1663_9.INJECT1_0 = "NO";
    defparam add_1663_9.INJECT1_1 = "NO";
    CCU2D add_1663_7 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [4]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [5]), 
          .D1(GND_net), .CIN(n27004), .COUT(n27005), .S0(n100[4]), .S1(n100[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_7.INIT0 = 16'h6969;
    defparam add_1663_7.INIT1 = 16'h6969;
    defparam add_1663_7.INJECT1_0 = "NO";
    defparam add_1663_7.INJECT1_1 = "NO";
    CCU2D add_1663_5 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [2]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [3]), 
          .D1(GND_net), .CIN(n27003), .COUT(n27004), .S0(n100[2]), .S1(n100[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_5.INIT0 = 16'h6969;
    defparam add_1663_5.INIT1 = 16'h6969;
    defparam add_1663_5.INJECT1_0 = "NO";
    defparam add_1663_5.INJECT1_1 = "NO";
    CCU2D add_1663_3 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [0]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [1]), 
          .D1(GND_net), .CIN(n27002), .COUT(n27003), .S0(n100[0]), .S1(n100[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_3.INIT0 = 16'h9696;
    defparam add_1663_3.INIT1 = 16'h6969;
    defparam add_1663_3.INJECT1_0 = "NO";
    defparam add_1663_3.INJECT1_1 = "NO";
    CCU2D add_1663_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(encoder_la_c), .B1(quadB_delayed), .C1(GND_net), .D1(GND_net), 
          .COUT(n27002));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_1.INIT0 = 16'hF000;
    defparam add_1663_1.INIT1 = 16'h6666;
    defparam add_1663_1.INJECT1_0 = "NO";
    defparam add_1663_1.INJECT1_1 = "NO";
    IFS1P3DX quadB_delayed_17 (.D(encoder_lb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam quadB_delayed_17.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_16 (.D(encoder_la_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam quadA_delayed_16.GSR = "ENABLED";
    CCU2D add_1663_33 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [30]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [31]), 
          .D1(GND_net), .CIN(n27017), .S0(n100[30]), .S1(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_33.INIT0 = 16'h6969;
    defparam add_1663_33.INIT1 = 16'h6969;
    defparam add_1663_33.INJECT1_0 = "NO";
    defparam add_1663_33.INJECT1_1 = "NO";
    CCU2D add_1663_31 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [28]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [29]), 
          .D1(GND_net), .CIN(n27016), .COUT(n27017), .S0(n100[28]), 
          .S1(n100[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_31.INIT0 = 16'h6969;
    defparam add_1663_31.INIT1 = 16'h6969;
    defparam add_1663_31.INJECT1_0 = "NO";
    defparam add_1663_31.INJECT1_1 = "NO";
    CCU2D add_1663_29 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [26]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [27]), 
          .D1(GND_net), .CIN(n27015), .COUT(n27016), .S0(n100[26]), 
          .S1(n100[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_29.INIT0 = 16'h6969;
    defparam add_1663_29.INIT1 = 16'h6969;
    defparam add_1663_29.INJECT1_0 = "NO";
    defparam add_1663_29.INJECT1_1 = "NO";
    LUT4 i14669_4_lut (.A(n31759), .B(encoder_la_c), .C(n6), .D(encoder_lb_c), 
         .Z(n13565)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i14669_4_lut.init = 16'hebbe;
    LUT4 i2_2_lut (.A(quadB_delayed), .B(quadA_delayed), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(17[22:59])
    defparam i2_2_lut.init = 16'h6666;
    CCU2D add_1663_27 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [24]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [25]), 
          .D1(GND_net), .CIN(n27014), .COUT(n27015), .S0(n100[24]), 
          .S1(n100[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_27.INIT0 = 16'h6969;
    defparam add_1663_27.INIT1 = 16'h6969;
    defparam add_1663_27.INJECT1_0 = "NO";
    defparam add_1663_27.INJECT1_1 = "NO";
    CCU2D add_1663_25 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [22]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [23]), 
          .D1(GND_net), .CIN(n27013), .COUT(n27014), .S0(n100[22]), 
          .S1(n100[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_25.INIT0 = 16'h6969;
    defparam add_1663_25.INIT1 = 16'h6969;
    defparam add_1663_25.INJECT1_0 = "NO";
    defparam add_1663_25.INJECT1_1 = "NO";
    CCU2D add_1663_23 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [20]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [21]), 
          .D1(GND_net), .CIN(n27012), .COUT(n27013), .S0(n100[20]), 
          .S1(n100[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_23.INIT0 = 16'h6969;
    defparam add_1663_23.INIT1 = 16'h6969;
    defparam add_1663_23.INJECT1_0 = "NO";
    defparam add_1663_23.INJECT1_1 = "NO";
    CCU2D add_1663_21 (.A0(encoder_la_c), .B0(quadB_delayed), .C0(\register[1] [18]), 
          .D0(GND_net), .A1(encoder_la_c), .B1(quadB_delayed), .C1(\register[1] [19]), 
          .D1(GND_net), .CIN(n27011), .COUT(n27012), .S0(n100[18]), 
          .S1(n100[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1663_21.INIT0 = 16'h6969;
    defparam add_1663_21.INIT1 = 16'h6969;
    defparam add_1663_21.INJECT1_0 = "NO";
    defparam add_1663_21.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module EncoderPeripheral
//

module EncoderPeripheral (n31780, n33457, \read_size[0] , n24748, encoder_ri_c, 
            \register_addr[0] , encoder_rb_c, encoder_ra_c, rw, n6, 
            n6_adj_14, n6_adj_15, n6_adj_16, n6_adj_17, n6_adj_18, 
            n6_adj_19, n6_adj_20, n6_adj_21, n6_adj_22, n6_adj_23, 
            n6_adj_24, n6_adj_25, n6_adj_26, n6_adj_27, n6_adj_28, 
            n6_adj_29, n6_adj_30, \read_value[1] , n31717, n31708, 
            \read_size[2] , n250, n8, n8_adj_31, n6_adj_32, n6_adj_33, 
            n6_adj_34, n6_adj_35, n6_adj_36, n6_adj_37, n8_adj_38, 
            n8_adj_39, n8_adj_40, n8_adj_41, n8_adj_42, debug_c_c, 
            n31759, n47, GND_net, n4144, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input n31780;
    input n33457;
    output \read_size[0] ;
    input n24748;
    input encoder_ri_c;
    input \register_addr[0] ;
    input encoder_rb_c;
    input encoder_ra_c;
    input rw;
    output n6;
    output n6_adj_14;
    output n6_adj_15;
    output n6_adj_16;
    output n6_adj_17;
    output n6_adj_18;
    output n6_adj_19;
    output n6_adj_20;
    output n6_adj_21;
    output n6_adj_22;
    output n6_adj_23;
    output n6_adj_24;
    output n6_adj_25;
    output n6_adj_26;
    output n6_adj_27;
    output n6_adj_28;
    output n6_adj_29;
    output n6_adj_30;
    output \read_value[1] ;
    input n31717;
    input n31708;
    output \read_size[2] ;
    input n250;
    output n8;
    output n8_adj_31;
    output n6_adj_32;
    output n6_adj_33;
    output n6_adj_34;
    output n6_adj_35;
    output n6_adj_36;
    output n6_adj_37;
    output n8_adj_38;
    output n8_adj_39;
    output n8_adj_40;
    output n8_adj_41;
    output n8_adj_42;
    input debug_c_c;
    input n31759;
    input n47;
    input GND_net;
    output n4144;
    input VCC_net;
    
    wire n31780 /* synthesis SET_AS_NETWORK=n31780 */ ;
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[13:23])
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(57[14:22])
    wire [31:0]n178;
    
    FD1S3IX read_value__i0 (.D(\register[1] [0]), .CK(n31780), .CD(n33457), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1S3AX read_size_i1 (.D(n24748), .CK(n31780), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 mux_113_Mux_1_i1_3_lut (.A(encoder_ri_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n178[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(76[29:42])
    defparam mux_113_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_113_Mux_2_i1_3_lut (.A(encoder_rb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n178[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(76[29:42])
    defparam mux_113_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_113_Mux_3_i1_3_lut (.A(encoder_ra_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n178[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(76[29:42])
    defparam mux_113_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 Select_4139_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[25]), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4139_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4157_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[19]), 
         .Z(n6_adj_14)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4157_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4142_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[24]), 
         .Z(n6_adj_15)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4142_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4145_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[23]), 
         .Z(n6_adj_16)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4145_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4148_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[22]), 
         .Z(n6_adj_17)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4148_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4151_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[21]), 
         .Z(n6_adj_18)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4151_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4154_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[20]), 
         .Z(n6_adj_19)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4154_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4160_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[18]), 
         .Z(n6_adj_20)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4160_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4163_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[17]), 
         .Z(n6_adj_21)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4163_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4166_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[16]), 
         .Z(n6_adj_22)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4166_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4169_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[15]), 
         .Z(n6_adj_23)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4169_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4172_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[14]), 
         .Z(n6_adj_24)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4172_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4175_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[13]), 
         .Z(n6_adj_25)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4175_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4178_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[12]), 
         .Z(n6_adj_26)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4178_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4181_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[11]), 
         .Z(n6_adj_27)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4181_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4184_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[10]), 
         .Z(n6_adj_28)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4184_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4187_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[9]), 
         .Z(n6_adj_29)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4187_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4190_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[8]), 
         .Z(n6_adj_30)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4190_i6_2_lut_3_lut.init = 16'h8080;
    FD1S3IX read_value__i1 (.D(n178[1]), .CK(n31780), .CD(n31717), .Q(\read_value[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n178[2]), .CK(n31780), .CD(n31717), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n178[3]), .CK(n31780), .CD(n31717), .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(\register[1] [4]), .CK(n31780), .CD(n33457), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(\register[1] [5]), .CK(n31780), .CD(n33457), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(\register[1] [6]), .CK(n31780), .CD(n33457), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i7 (.D(\register[1] [7]), .CK(n31780), .CD(n33457), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1S3IX read_value__i8 (.D(\register[1] [8]), .CK(n31780), .CD(n33457), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1S3IX read_value__i9 (.D(\register[1] [9]), .CK(n31780), .CD(n33457), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1S3IX read_value__i10 (.D(\register[1] [10]), .CK(n31780), .CD(n33457), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1S3IX read_value__i11 (.D(\register[1] [11]), .CK(n31780), .CD(n33457), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1S3IX read_value__i12 (.D(\register[1] [12]), .CK(n31780), .CD(n33457), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1S3IX read_value__i13 (.D(\register[1] [13]), .CK(n31780), .CD(n33457), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1S3IX read_value__i14 (.D(\register[1] [14]), .CK(n31780), .CD(n33457), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1S3IX read_value__i15 (.D(\register[1] [15]), .CK(n31780), .CD(n33457), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1S3IX read_value__i16 (.D(\register[1] [16]), .CK(n31780), .CD(n33457), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1S3IX read_value__i17 (.D(\register[1] [17]), .CK(n31780), .CD(n33457), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1S3IX read_value__i18 (.D(\register[1] [18]), .CK(n31780), .CD(n33457), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1S3IX read_value__i19 (.D(\register[1] [19]), .CK(n31780), .CD(n33457), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1S3IX read_value__i20 (.D(\register[1] [20]), .CK(n31780), .CD(n33457), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1S3IX read_value__i21 (.D(\register[1] [21]), .CK(n31780), .CD(n33457), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1S3IX read_value__i22 (.D(\register[1] [22]), .CK(n31780), .CD(n33457), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1S3IX read_value__i23 (.D(\register[1] [23]), .CK(n31780), .CD(n33457), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1S3IX read_value__i24 (.D(\register[1] [24]), .CK(n31780), .CD(n31708), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1S3IX read_value__i25 (.D(\register[1] [25]), .CK(n31780), .CD(n31708), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1S3IX read_value__i26 (.D(\register[1] [26]), .CK(n31780), .CD(n31708), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1S3IX read_value__i27 (.D(\register[1] [27]), .CK(n31780), .CD(n31708), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1S3IX read_value__i28 (.D(\register[1] [28]), .CK(n31780), .CD(n31708), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1S3IX read_value__i29 (.D(\register[1] [29]), .CK(n31780), .CD(n31708), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1S3IX read_value__i30 (.D(\register[1] [30]), .CK(n31780), .CD(n31708), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1S3IX read_value__i31 (.D(\register[1] [31]), .CK(n31780), .CD(n31708), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1S3AX read_size_i2 (.D(n250), .CK(n31780), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=657, LSE_RLINE=667 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 84[6])
    defparam read_size_i2.GSR = "ENABLED";
    LUT4 Select_4196_i8_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[2]), 
         .Z(n8)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4196_i8_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4198_i8_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[0]), 
         .Z(n8_adj_31)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4198_i8_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4121_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[31]), 
         .Z(n6_adj_32)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4121_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4124_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[30]), 
         .Z(n6_adj_33)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4124_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4127_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[29]), 
         .Z(n6_adj_34)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4127_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4130_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[28]), 
         .Z(n6_adj_35)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4130_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4133_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[27]), 
         .Z(n6_adj_36)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4133_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4136_i6_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[26]), 
         .Z(n6_adj_37)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4136_i6_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4191_i8_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[7]), 
         .Z(n8_adj_38)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4191_i8_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4192_i8_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[6]), 
         .Z(n8_adj_39)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4192_i8_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4193_i8_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[5]), 
         .Z(n8_adj_40)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4193_i8_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4194_i8_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[4]), 
         .Z(n8_adj_41)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4194_i8_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4195_i8_2_lut_3_lut (.A(n31780), .B(rw), .C(read_value[3]), 
         .Z(n8_adj_42)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(69[19:32])
    defparam Select_4195_i8_2_lut_3_lut.init = 16'h8080;
    QuadratureDecoder q (.\register[1] ({\register[1] }), .debug_c_c(debug_c_c), 
            .n31759(n31759), .n47(n47), .encoder_ra_c(encoder_ra_c), .GND_net(GND_net), 
            .n4144(n4144), .encoder_rb_c(encoder_rb_c), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(88[20] 92[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder
//

module QuadratureDecoder (\register[1] , debug_c_c, n31759, n47, encoder_ra_c, 
            GND_net, n4144, encoder_rb_c, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[1] ;
    input debug_c_c;
    input n31759;
    input n47;
    input encoder_ra_c;
    input GND_net;
    output n4144;
    input encoder_rb_c;
    input VCC_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n13611;
    wire [31:0]n100;
    
    wire n27684, quadB_delayed, n27683, n27682, n27681, n27680, 
        n27679, n27678, n6, quadA_delayed, n27677, n27676, n27675, 
        n27674, n27673, n27672, n27671, n27670, n27669;
    
    FD1P3IX count__i21 (.D(n100[21]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i31 (.D(n100[31]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n100[30]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n100[29]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n100[28]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n100[27]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n100[26]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3AX count__i25 (.D(n47), .SP(n13611), .CK(debug_c_c), .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n100[24]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n100[23]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n100[22]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n100[20]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n100[19]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n100[18]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n100[17]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n100[16]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n100[15]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n100[14]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n100[13]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n100[12]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n100[11]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n100[10]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n100[9]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n100[8]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n100[7]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n100[6]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n100[5]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n100[4]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n100[3]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n100[2]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n100[1]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i0 (.D(n100[0]), .SP(n13611), .CD(n31759), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_1629_33 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [30]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [31]), 
          .D1(GND_net), .CIN(n27684), .S0(n100[30]), .S1(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_33.INIT0 = 16'h6969;
    defparam add_1629_33.INIT1 = 16'h6969;
    defparam add_1629_33.INJECT1_0 = "NO";
    defparam add_1629_33.INJECT1_1 = "NO";
    CCU2D add_1629_31 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [28]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [29]), 
          .D1(GND_net), .CIN(n27683), .COUT(n27684), .S0(n100[28]), 
          .S1(n100[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_31.INIT0 = 16'h6969;
    defparam add_1629_31.INIT1 = 16'h6969;
    defparam add_1629_31.INJECT1_0 = "NO";
    defparam add_1629_31.INJECT1_1 = "NO";
    CCU2D add_1629_29 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [26]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [27]), 
          .D1(GND_net), .CIN(n27682), .COUT(n27683), .S0(n100[26]), 
          .S1(n100[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_29.INIT0 = 16'h6969;
    defparam add_1629_29.INIT1 = 16'h6969;
    defparam add_1629_29.INJECT1_0 = "NO";
    defparam add_1629_29.INJECT1_1 = "NO";
    CCU2D add_1629_27 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [24]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [25]), 
          .D1(GND_net), .CIN(n27681), .COUT(n27682), .S0(n100[24]), 
          .S1(n4144));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_27.INIT0 = 16'h6969;
    defparam add_1629_27.INIT1 = 16'h6969;
    defparam add_1629_27.INJECT1_0 = "NO";
    defparam add_1629_27.INJECT1_1 = "NO";
    CCU2D add_1629_25 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [22]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [23]), 
          .D1(GND_net), .CIN(n27680), .COUT(n27681), .S0(n100[22]), 
          .S1(n100[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_25.INIT0 = 16'h6969;
    defparam add_1629_25.INIT1 = 16'h6969;
    defparam add_1629_25.INJECT1_0 = "NO";
    defparam add_1629_25.INJECT1_1 = "NO";
    CCU2D add_1629_23 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [20]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [21]), 
          .D1(GND_net), .CIN(n27679), .COUT(n27680), .S0(n100[20]), 
          .S1(n100[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_23.INIT0 = 16'h6969;
    defparam add_1629_23.INIT1 = 16'h6969;
    defparam add_1629_23.INJECT1_0 = "NO";
    defparam add_1629_23.INJECT1_1 = "NO";
    CCU2D add_1629_21 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [18]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [19]), 
          .D1(GND_net), .CIN(n27678), .COUT(n27679), .S0(n100[18]), 
          .S1(n100[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_21.INIT0 = 16'h6969;
    defparam add_1629_21.INIT1 = 16'h6969;
    defparam add_1629_21.INJECT1_0 = "NO";
    defparam add_1629_21.INJECT1_1 = "NO";
    LUT4 i14667_4_lut (.A(n31759), .B(encoder_ra_c), .C(n6), .D(encoder_rb_c), 
         .Z(n13611)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i14667_4_lut.init = 16'hebbe;
    LUT4 i2_2_lut (.A(quadB_delayed), .B(quadA_delayed), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(17[22:59])
    defparam i2_2_lut.init = 16'h6666;
    IFS1P3DX quadB_delayed_17 (.D(encoder_rb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam quadB_delayed_17.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_16 (.D(encoder_ra_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=88, LSE_RLINE=92 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 36[6])
    defparam quadA_delayed_16.GSR = "ENABLED";
    CCU2D add_1629_19 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [16]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [17]), 
          .D1(GND_net), .CIN(n27677), .COUT(n27678), .S0(n100[16]), 
          .S1(n100[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_19.INIT0 = 16'h6969;
    defparam add_1629_19.INIT1 = 16'h6969;
    defparam add_1629_19.INJECT1_0 = "NO";
    defparam add_1629_19.INJECT1_1 = "NO";
    CCU2D add_1629_17 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [14]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [15]), 
          .D1(GND_net), .CIN(n27676), .COUT(n27677), .S0(n100[14]), 
          .S1(n100[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_17.INIT0 = 16'h6969;
    defparam add_1629_17.INIT1 = 16'h6969;
    defparam add_1629_17.INJECT1_0 = "NO";
    defparam add_1629_17.INJECT1_1 = "NO";
    CCU2D add_1629_15 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [12]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [13]), 
          .D1(GND_net), .CIN(n27675), .COUT(n27676), .S0(n100[12]), 
          .S1(n100[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_15.INIT0 = 16'h6969;
    defparam add_1629_15.INIT1 = 16'h6969;
    defparam add_1629_15.INJECT1_0 = "NO";
    defparam add_1629_15.INJECT1_1 = "NO";
    CCU2D add_1629_13 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [10]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [11]), 
          .D1(GND_net), .CIN(n27674), .COUT(n27675), .S0(n100[10]), 
          .S1(n100[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_13.INIT0 = 16'h6969;
    defparam add_1629_13.INIT1 = 16'h6969;
    defparam add_1629_13.INJECT1_0 = "NO";
    defparam add_1629_13.INJECT1_1 = "NO";
    CCU2D add_1629_11 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [8]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [9]), 
          .D1(GND_net), .CIN(n27673), .COUT(n27674), .S0(n100[8]), .S1(n100[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_11.INIT0 = 16'h6969;
    defparam add_1629_11.INIT1 = 16'h6969;
    defparam add_1629_11.INJECT1_0 = "NO";
    defparam add_1629_11.INJECT1_1 = "NO";
    CCU2D add_1629_9 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [6]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [7]), 
          .D1(GND_net), .CIN(n27672), .COUT(n27673), .S0(n100[6]), .S1(n100[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_9.INIT0 = 16'h6969;
    defparam add_1629_9.INIT1 = 16'h6969;
    defparam add_1629_9.INJECT1_0 = "NO";
    defparam add_1629_9.INJECT1_1 = "NO";
    CCU2D add_1629_7 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [4]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [5]), 
          .D1(GND_net), .CIN(n27671), .COUT(n27672), .S0(n100[4]), .S1(n100[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_7.INIT0 = 16'h6969;
    defparam add_1629_7.INIT1 = 16'h6969;
    defparam add_1629_7.INJECT1_0 = "NO";
    defparam add_1629_7.INJECT1_1 = "NO";
    CCU2D add_1629_5 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [2]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [3]), 
          .D1(GND_net), .CIN(n27670), .COUT(n27671), .S0(n100[2]), .S1(n100[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_5.INIT0 = 16'h6969;
    defparam add_1629_5.INIT1 = 16'h6969;
    defparam add_1629_5.INJECT1_0 = "NO";
    defparam add_1629_5.INJECT1_1 = "NO";
    CCU2D add_1629_3 (.A0(encoder_ra_c), .B0(quadB_delayed), .C0(\register[1] [0]), 
          .D0(GND_net), .A1(encoder_ra_c), .B1(quadB_delayed), .C1(\register[1] [1]), 
          .D1(GND_net), .CIN(n27669), .COUT(n27670), .S0(n100[0]), .S1(n100[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_3.INIT0 = 16'h9696;
    defparam add_1629_3.INIT1 = 16'h6969;
    defparam add_1629_3.INJECT1_0 = "NO";
    defparam add_1629_3.INJECT1_1 = "NO";
    CCU2D add_1629_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(encoder_ra_c), .B1(quadB_delayed), .C1(GND_net), .D1(GND_net), 
          .COUT(n27669));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(30[5] 35[8])
    defparam add_1629_1.INIT0 = 16'hF000;
    defparam add_1629_1.INIT1 = 16'h6666;
    defparam add_1629_1.INJECT1_0 = "NO";
    defparam add_1629_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (GND_net, debug_c_c, VCC_net, 
            Stepper_Y_nFault_c, n33450, \read_size[0] , n14194, n78, 
            Stepper_Y_M0_c_0, n89, n579, prev_step_clk, step_clk, 
            n14084, prev_select, n31727, \steps_reg[9] , \steps_reg[5] , 
            \steps_reg[6] , \steps_reg[3] , n32, \register_addr[0] , 
            n27893, Stepper_Y_M1_c_1, int_step, n22, n31712, n31724, 
            n33448, databus, n33451, n33452, \div_factor_reg[9] , 
            \div_factor_reg[6] , \div_factor_reg[5] , \div_factor_reg[3] , 
            \control_reg[7] , n13606, Stepper_Y_En_c, Stepper_Y_Dir_c, 
            \control_reg[3] , Stepper_Y_M2_c_2, \read_size[2] , n33453, 
            read_value, \register_addr[1] , n8243, n3883, n33447, 
            limit_c_1, n31785, \register_addr[3] , \register_addr[2] , 
            n79, n6584, n20993, n20982) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input VCC_net;
    input Stepper_Y_nFault_c;
    input n33450;
    output \read_size[0] ;
    input n14194;
    input n78;
    output Stepper_Y_M0_c_0;
    input n89;
    input n579;
    output prev_step_clk;
    output step_clk;
    input n14084;
    output prev_select;
    input n31727;
    output \steps_reg[9] ;
    output \steps_reg[5] ;
    output \steps_reg[6] ;
    output \steps_reg[3] ;
    input n32;
    input \register_addr[0] ;
    output n27893;
    output Stepper_Y_M1_c_1;
    output int_step;
    input n22;
    input n31712;
    input n31724;
    input n33448;
    input [31:0]databus;
    input n33451;
    input n33452;
    output \div_factor_reg[9] ;
    output \div_factor_reg[6] ;
    output \div_factor_reg[5] ;
    output \div_factor_reg[3] ;
    output \control_reg[7] ;
    input n13606;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output \control_reg[3] ;
    output Stepper_Y_M2_c_2;
    output \read_size[2] ;
    input n33453;
    output [31:0]read_value;
    input \register_addr[1] ;
    input n8243;
    input n3883;
    input n33447;
    input limit_c_1;
    input n31785;
    input \register_addr[3] ;
    input \register_addr[2] ;
    input n79;
    input n6584;
    input n20993;
    input n20982;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27362;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n224;
    
    wire n27361, fault_latched;
    wire [31:0]n3884;
    
    wire limit_latched, n182, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n27360, n27359, n27358, n27357, n27356, n27355, n27354, 
        n27353, n27352, n27351, n27350, n27349, n27348, n27347, 
        n30080, n30081, n49, n62, n58, n50, n41, n60, n54, 
        n42, n52, n38, n56, n46, n30101, n30102, n11642;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n27972, n30050, n30051, n30052;
    wire [7:0]n8242;
    wire [31:0]n6522;
    wire [31:0]n6558;
    wire [31:0]n99;
    
    wire n30082, n30103;
    
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27362), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27361), .COUT(n27362), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3884[0]), .CK(debug_c_c), .CD(n33450), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n78), .SP(n14194), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n89), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n14084), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31727), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27360), .COUT(n27361), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27359), .COUT(n27360), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27358), .COUT(n27359), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27357), .COUT(n27358), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27356), .COUT(n27357), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27355), .COUT(n27356), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27354), .COUT(n27355), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27353), .COUT(n27354), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27352), .COUT(n27353), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27351), .COUT(n27352), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27350), .COUT(n27351), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27349), .COUT(n27350), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27348), .COUT(n27349), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27347), .COUT(n27348), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27347), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i22927_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22927_3_lut.init = 16'hcaca;
    LUT4 i22928_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22928_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27893)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22948_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22948_3_lut.init = 16'hcaca;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i22949_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22949_3_lut.init = 16'hcaca;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    FD1P3AX int_step_182 (.D(n31712), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n31724), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n31724), .CD(n33451), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n31724), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n31724), .CD(n33451), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n31724), .PD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n31724), .PD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n31724), .PD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n31724), .PD(n33452), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n31724), .PD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n31724), .PD(n33448), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n31724), .PD(n33448), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n31724), .CD(n33452), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n31724), .CD(n33448), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n31724), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n31724), .CD(n33448), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13606), .CD(n11642), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13606), .PD(n33448), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13606), .PD(n33452), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13606), .CD(n33452), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13606), .PD(n33448), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13606), .CD(n33448), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13606), .PD(n33448), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n27972), .SP(n14194), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3884[31]), .CK(debug_c_c), .CD(n33448), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3884[30]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3884[29]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3884[28]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3884[27]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3884[26]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3884[25]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3884[24]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3884[23]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3884[22]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3884[21]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3884[20]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3884[19]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3884[18]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3884[17]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3884[16]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3884[15]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3884[14]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3884[13]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3884[12]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3884[11]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3884[10]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3884[9]), .CK(debug_c_c), .CD(n33452), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3884[8]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3884[7]), .CK(debug_c_c), .CD(n33452), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3884[6]), .CK(debug_c_c), .CD(n33453), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3884[5]), .CK(debug_c_c), .CD(n33453), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3884[4]), .CK(debug_c_c), .CD(n33453), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3884[3]), .CK(debug_c_c), .CD(n33453), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3884[2]), .CK(debug_c_c), .CD(n33453), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3884[1]), .CK(debug_c_c), .CD(n33453), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    PFUMX i22899 (.BLUT(n30050), .ALUT(n30051), .C0(\register_addr[0] ), 
          .Z(n30052));
    LUT4 i14864_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8242[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14864_2_lut.init = 16'h2222;
    LUT4 mux_1895_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n6522[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1895_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1895_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6522[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1895_i8_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i11 (.D(n6558[11]), .SP(n14194), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n6558[12]), .SP(n14194), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n6558[13]), .SP(n14194), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n6558[14]), .SP(n14194), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n6558[15]), .SP(n14194), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n6558[16]), .SP(n14194), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n6558[17]), .SP(n14194), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    LUT4 i14995_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n99[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14995_4_lut.init = 16'hc088;
    LUT4 i14992_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n99[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14992_4_lut.init = 16'hc088;
    LUT4 i14991_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n99[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14991_4_lut.init = 16'hc088;
    LUT4 i14990_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n99[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14990_4_lut.init = 16'hc088;
    LUT4 i14989_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n99[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14989_4_lut.init = 16'hc088;
    LUT4 i14988_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n99[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14988_4_lut.init = 16'hc088;
    LUT4 i14985_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n99[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14985_4_lut.init = 16'hc088;
    LUT4 i15178_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n99[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15178_4_lut.init = 16'hc088;
    LUT4 i15177_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n99[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15177_4_lut.init = 16'hc088;
    LUT4 i14998_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n99[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14998_4_lut.init = 16'hc088;
    LUT4 i15176_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n99[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15176_4_lut.init = 16'hc088;
    LUT4 i15175_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n99[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15175_4_lut.init = 16'hc088;
    LUT4 i15174_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n99[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15174_4_lut.init = 16'hc088;
    LUT4 i15173_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n99[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15173_4_lut.init = 16'hc088;
    LUT4 i14954_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n99[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14954_4_lut.init = 16'hc088;
    LUT4 i14949_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n99[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i14949_4_lut.init = 16'hc088;
    PFUMX i22929 (.BLUT(n30080), .ALUT(n30081), .C0(\register_addr[1] ), 
          .Z(n30082));
    PFUMX i22950 (.BLUT(n30101), .ALUT(n30102), .C0(\register_addr[1] ), 
          .Z(n30103));
    PFUMX mux_1899_i5 (.BLUT(n8242[4]), .ALUT(n6522[4]), .C0(\register_addr[1] ), 
          .Z(n6558[4]));
    PFUMX mux_1899_i8 (.BLUT(n8243), .ALUT(n6522[7]), .C0(\register_addr[1] ), 
          .Z(n6558[7]));
    LUT4 mux_1546_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3883), .Z(n3884[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n30082), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30103), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30052), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n99[31]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n99[30]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n99[29]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n99[28]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n99[27]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n99[26]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n99[25]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n99[24]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    LUT4 i22897_3_lut (.A(Stepper_Y_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22897_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i23 (.D(n99[23]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n99[22]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    LUT4 i5242_3_lut (.A(prev_limit_latched), .B(n33447), .C(limit_latched), 
         .Z(n11642)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i5242_3_lut.init = 16'hdcdc;
    LUT4 i22898_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22898_3_lut.init = 16'hcaca;
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i23093_4_lut (.A(n31785), .B(\register_addr[1] ), .C(\register_addr[3] ), 
         .D(\register_addr[2] ), .Z(n27972)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i23093_4_lut.init = 16'h0004;
    LUT4 mux_1546_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3883), 
         .Z(n3884[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3883), 
         .Z(n3884[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3883), 
         .Z(n3884[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3883), 
         .Z(n3884[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3883), 
         .Z(n3884[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3883), 
         .Z(n3884[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3883), 
         .Z(n3884[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3883), 
         .Z(n3884[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3883), 
         .Z(n3884[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3883), 
         .Z(n3884[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3883), 
         .Z(n3884[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3883), 
         .Z(n3884[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3883), 
         .Z(n3884[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3883), 
         .Z(n3884[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3883), 
         .Z(n3884[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3883), 
         .Z(n3884[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3883), 
         .Z(n3884[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3883), 
         .Z(n3884[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3883), 
         .Z(n3884[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3883), 
         .Z(n3884[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3883), 
         .Z(n3884[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3883), 
         .Z(n3884[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3883), .Z(n3884[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3883), .Z(n3884[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3883), .Z(n3884[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3883), .Z(n3884[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3883), .Z(n3884[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3883), .Z(n3884[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3883), .Z(n3884[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3883), .Z(n3884[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1546_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3883), .Z(n3884[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1546_i2_3_lut.init = 16'hcaca;
    LUT4 i14871_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n6558[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14871_4_lut.init = 16'hc088;
    LUT4 i14870_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n6558[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14870_4_lut.init = 16'hc088;
    LUT4 i14869_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n6558[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14869_4_lut.init = 16'hc088;
    LUT4 i14868_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n6558[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14868_4_lut.init = 16'hc088;
    LUT4 i14867_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n6558[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14867_4_lut.init = 16'hc088;
    LUT4 i14866_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n6558[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14866_4_lut.init = 16'hc088;
    LUT4 i14865_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n6558[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14865_4_lut.init = 16'hc088;
    FD1P3AX read_value__i21 (.D(n99[21]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n99[20]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n99[19]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n99[18]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n99[10]), .SP(n14194), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n79), .SP(n14194), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n99[8]), .SP(n14194), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6558[7]), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6584), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n20993), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6558[4]), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n20982), .SP(n14194), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=573, LSE_RLINE=586 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    ClockDivider_U7 step_clk_gen (.n33447(n33447), .debug_c_c(debug_c_c), 
            .div_factor_reg({div_factor_reg[31:10], \div_factor_reg[9] , 
            div_factor_reg[8:7], \div_factor_reg[6] , \div_factor_reg[5] , 
            div_factor_reg[4], \div_factor_reg[3] , div_factor_reg[2:0]}), 
            .GND_net(GND_net), .step_clk(step_clk), .n33448(n33448)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (n33447, debug_c_c, div_factor_reg, GND_net, 
            step_clk, n33448) /* synthesis syn_module_defined=1 */ ;
    input n33447;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input GND_net;
    output step_clk;
    input n33448;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7763, n31693;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n16110, n27162;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n7728, n27161, n27160, n27159, n27158, n27157, n27156, 
        n27155, n27154, n27153, n27152, n27151, n27150, n27149, 
        n27148, n27147, n27146;
    wire [31:0]n40;
    
    wire n27145, n27144, n27143, n27142, n27141, n27140, n27139, 
        n27138, n27137, n27136, n27135, n27134, n27133, n7797, 
        n27132, n27131, n27130, n27129, n27128, n27127;
    wire [31:0]n134;
    
    wire n27126, n27125, n27124, n27123, n27122, n27121, n27120, 
        n27119, n27118, n27117, n27116, n27115, n27298, n27297, 
        n27296, n27295, n27294, n27293, n27292, n27291, n27290, 
        n27289, n27288, n27287, n27402, n27286, n27285, n27401, 
        n27284, n27400, n27399, n27398, n27283, n27397, n27396, 
        n27395, n27394, n27393, n27392, n27391, n27390, n27389, 
        n27388, n27387;
    
    LUT4 i1005_2_lut_rep_270 (.A(n7763), .B(n33447), .Z(n31693)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1005_2_lut_rep_270.init = 16'heeee;
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_1999_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27162), .S1(n7728));
    defparam sub_1999_add_2_33.INIT0 = 16'h5555;
    defparam sub_1999_add_2_33.INIT1 = 16'h0000;
    defparam sub_1999_add_2_33.INJECT1_0 = "NO";
    defparam sub_1999_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27161), .COUT(n27162));
    defparam sub_1999_add_2_31.INIT0 = 16'h5999;
    defparam sub_1999_add_2_31.INIT1 = 16'h5999;
    defparam sub_1999_add_2_31.INJECT1_0 = "NO";
    defparam sub_1999_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27160), .COUT(n27161));
    defparam sub_1999_add_2_29.INIT0 = 16'h5999;
    defparam sub_1999_add_2_29.INIT1 = 16'h5999;
    defparam sub_1999_add_2_29.INJECT1_0 = "NO";
    defparam sub_1999_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27159), .COUT(n27160));
    defparam sub_1999_add_2_27.INIT0 = 16'h5999;
    defparam sub_1999_add_2_27.INIT1 = 16'h5999;
    defparam sub_1999_add_2_27.INJECT1_0 = "NO";
    defparam sub_1999_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27158), .COUT(n27159));
    defparam sub_1999_add_2_25.INIT0 = 16'h5999;
    defparam sub_1999_add_2_25.INIT1 = 16'h5999;
    defparam sub_1999_add_2_25.INJECT1_0 = "NO";
    defparam sub_1999_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27157), .COUT(n27158));
    defparam sub_1999_add_2_23.INIT0 = 16'h5999;
    defparam sub_1999_add_2_23.INIT1 = 16'h5999;
    defparam sub_1999_add_2_23.INJECT1_0 = "NO";
    defparam sub_1999_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27156), .COUT(n27157));
    defparam sub_1999_add_2_21.INIT0 = 16'h5999;
    defparam sub_1999_add_2_21.INIT1 = 16'h5999;
    defparam sub_1999_add_2_21.INJECT1_0 = "NO";
    defparam sub_1999_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27155), .COUT(n27156));
    defparam sub_1999_add_2_19.INIT0 = 16'h5999;
    defparam sub_1999_add_2_19.INIT1 = 16'h5999;
    defparam sub_1999_add_2_19.INJECT1_0 = "NO";
    defparam sub_1999_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27154), .COUT(n27155));
    defparam sub_1999_add_2_17.INIT0 = 16'h5999;
    defparam sub_1999_add_2_17.INIT1 = 16'h5999;
    defparam sub_1999_add_2_17.INJECT1_0 = "NO";
    defparam sub_1999_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27153), .COUT(n27154));
    defparam sub_1999_add_2_15.INIT0 = 16'h5999;
    defparam sub_1999_add_2_15.INIT1 = 16'h5999;
    defparam sub_1999_add_2_15.INJECT1_0 = "NO";
    defparam sub_1999_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27152), .COUT(n27153));
    defparam sub_1999_add_2_13.INIT0 = 16'h5999;
    defparam sub_1999_add_2_13.INIT1 = 16'h5999;
    defparam sub_1999_add_2_13.INJECT1_0 = "NO";
    defparam sub_1999_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27151), .COUT(n27152));
    defparam sub_1999_add_2_11.INIT0 = 16'h5999;
    defparam sub_1999_add_2_11.INIT1 = 16'h5999;
    defparam sub_1999_add_2_11.INJECT1_0 = "NO";
    defparam sub_1999_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27150), .COUT(n27151));
    defparam sub_1999_add_2_9.INIT0 = 16'h5999;
    defparam sub_1999_add_2_9.INIT1 = 16'h5999;
    defparam sub_1999_add_2_9.INJECT1_0 = "NO";
    defparam sub_1999_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27149), .COUT(n27150));
    defparam sub_1999_add_2_7.INIT0 = 16'h5999;
    defparam sub_1999_add_2_7.INIT1 = 16'h5999;
    defparam sub_1999_add_2_7.INJECT1_0 = "NO";
    defparam sub_1999_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27148), .COUT(n27149));
    defparam sub_1999_add_2_5.INIT0 = 16'h5999;
    defparam sub_1999_add_2_5.INIT1 = 16'h5999;
    defparam sub_1999_add_2_5.INJECT1_0 = "NO";
    defparam sub_1999_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27147), .COUT(n27148));
    defparam sub_1999_add_2_3.INIT0 = 16'h5999;
    defparam sub_1999_add_2_3.INIT1 = 16'h5999;
    defparam sub_1999_add_2_3.INJECT1_0 = "NO";
    defparam sub_1999_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1999_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27147));
    defparam sub_1999_add_2_1.INIT0 = 16'h0000;
    defparam sub_1999_add_2_1.INIT1 = 16'h5999;
    defparam sub_1999_add_2_1.INJECT1_0 = "NO";
    defparam sub_1999_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27146), .S1(n7763));
    defparam sub_2001_add_2_33.INIT0 = 16'h5999;
    defparam sub_2001_add_2_33.INIT1 = 16'h0000;
    defparam sub_2001_add_2_33.INJECT1_0 = "NO";
    defparam sub_2001_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27145), .COUT(n27146));
    defparam sub_2001_add_2_31.INIT0 = 16'h5999;
    defparam sub_2001_add_2_31.INIT1 = 16'h5999;
    defparam sub_2001_add_2_31.INJECT1_0 = "NO";
    defparam sub_2001_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27144), .COUT(n27145));
    defparam sub_2001_add_2_29.INIT0 = 16'h5999;
    defparam sub_2001_add_2_29.INIT1 = 16'h5999;
    defparam sub_2001_add_2_29.INJECT1_0 = "NO";
    defparam sub_2001_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27143), .COUT(n27144));
    defparam sub_2001_add_2_27.INIT0 = 16'h5999;
    defparam sub_2001_add_2_27.INIT1 = 16'h5999;
    defparam sub_2001_add_2_27.INJECT1_0 = "NO";
    defparam sub_2001_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27142), .COUT(n27143));
    defparam sub_2001_add_2_25.INIT0 = 16'h5999;
    defparam sub_2001_add_2_25.INIT1 = 16'h5999;
    defparam sub_2001_add_2_25.INJECT1_0 = "NO";
    defparam sub_2001_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27141), .COUT(n27142));
    defparam sub_2001_add_2_23.INIT0 = 16'h5999;
    defparam sub_2001_add_2_23.INIT1 = 16'h5999;
    defparam sub_2001_add_2_23.INJECT1_0 = "NO";
    defparam sub_2001_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27140), .COUT(n27141));
    defparam sub_2001_add_2_21.INIT0 = 16'h5999;
    defparam sub_2001_add_2_21.INIT1 = 16'h5999;
    defparam sub_2001_add_2_21.INJECT1_0 = "NO";
    defparam sub_2001_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27139), .COUT(n27140));
    defparam sub_2001_add_2_19.INIT0 = 16'h5999;
    defparam sub_2001_add_2_19.INIT1 = 16'h5999;
    defparam sub_2001_add_2_19.INJECT1_0 = "NO";
    defparam sub_2001_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27138), .COUT(n27139));
    defparam sub_2001_add_2_17.INIT0 = 16'h5999;
    defparam sub_2001_add_2_17.INIT1 = 16'h5999;
    defparam sub_2001_add_2_17.INJECT1_0 = "NO";
    defparam sub_2001_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27137), .COUT(n27138));
    defparam sub_2001_add_2_15.INIT0 = 16'h5999;
    defparam sub_2001_add_2_15.INIT1 = 16'h5999;
    defparam sub_2001_add_2_15.INJECT1_0 = "NO";
    defparam sub_2001_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27136), .COUT(n27137));
    defparam sub_2001_add_2_13.INIT0 = 16'h5999;
    defparam sub_2001_add_2_13.INIT1 = 16'h5999;
    defparam sub_2001_add_2_13.INJECT1_0 = "NO";
    defparam sub_2001_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27135), .COUT(n27136));
    defparam sub_2001_add_2_11.INIT0 = 16'h5999;
    defparam sub_2001_add_2_11.INIT1 = 16'h5999;
    defparam sub_2001_add_2_11.INJECT1_0 = "NO";
    defparam sub_2001_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27134), .COUT(n27135));
    defparam sub_2001_add_2_9.INIT0 = 16'h5999;
    defparam sub_2001_add_2_9.INIT1 = 16'h5999;
    defparam sub_2001_add_2_9.INJECT1_0 = "NO";
    defparam sub_2001_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27133), .COUT(n27134));
    defparam sub_2001_add_2_7.INIT0 = 16'h5999;
    defparam sub_2001_add_2_7.INIT1 = 16'h5999;
    defparam sub_2001_add_2_7.INJECT1_0 = "NO";
    defparam sub_2001_add_2_7.INJECT1_1 = "NO";
    LUT4 i9704_2_lut_3_lut (.A(n7763), .B(n33447), .C(n7797), .Z(n16110)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i9704_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_2001_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27132), .COUT(n27133));
    defparam sub_2001_add_2_5.INIT0 = 16'h5999;
    defparam sub_2001_add_2_5.INIT1 = 16'h5999;
    defparam sub_2001_add_2_5.INJECT1_0 = "NO";
    defparam sub_2001_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27131), .COUT(n27132));
    defparam sub_2001_add_2_3.INIT0 = 16'h5999;
    defparam sub_2001_add_2_3.INIT1 = 16'h5999;
    defparam sub_2001_add_2_3.INJECT1_0 = "NO";
    defparam sub_2001_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2001_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27131));
    defparam sub_2001_add_2_1.INIT0 = 16'h0000;
    defparam sub_2001_add_2_1.INIT1 = 16'h5999;
    defparam sub_2001_add_2_1.INJECT1_0 = "NO";
    defparam sub_2001_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27130), .S1(n7797));
    defparam sub_2002_add_2_33.INIT0 = 16'hf555;
    defparam sub_2002_add_2_33.INIT1 = 16'h0000;
    defparam sub_2002_add_2_33.INJECT1_0 = "NO";
    defparam sub_2002_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27129), .COUT(n27130));
    defparam sub_2002_add_2_31.INIT0 = 16'hf555;
    defparam sub_2002_add_2_31.INIT1 = 16'hf555;
    defparam sub_2002_add_2_31.INJECT1_0 = "NO";
    defparam sub_2002_add_2_31.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7728), .CK(debug_c_c), .CD(n33448), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2002_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27128), .COUT(n27129));
    defparam sub_2002_add_2_29.INIT0 = 16'hf555;
    defparam sub_2002_add_2_29.INIT1 = 16'hf555;
    defparam sub_2002_add_2_29.INJECT1_0 = "NO";
    defparam sub_2002_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27127), .COUT(n27128));
    defparam sub_2002_add_2_27.INIT0 = 16'hf555;
    defparam sub_2002_add_2_27.INIT1 = 16'hf555;
    defparam sub_2002_add_2_27.INJECT1_0 = "NO";
    defparam sub_2002_add_2_27.INJECT1_1 = "NO";
    FD1S3IX count_2579__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i0.GSR = "ENABLED";
    CCU2D sub_2002_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27126), .COUT(n27127));
    defparam sub_2002_add_2_25.INIT0 = 16'hf555;
    defparam sub_2002_add_2_25.INIT1 = 16'hf555;
    defparam sub_2002_add_2_25.INJECT1_0 = "NO";
    defparam sub_2002_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27125), .COUT(n27126));
    defparam sub_2002_add_2_23.INIT0 = 16'hf555;
    defparam sub_2002_add_2_23.INIT1 = 16'hf555;
    defparam sub_2002_add_2_23.INJECT1_0 = "NO";
    defparam sub_2002_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27124), .COUT(n27125));
    defparam sub_2002_add_2_21.INIT0 = 16'hf555;
    defparam sub_2002_add_2_21.INIT1 = 16'hf555;
    defparam sub_2002_add_2_21.INJECT1_0 = "NO";
    defparam sub_2002_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27123), .COUT(n27124));
    defparam sub_2002_add_2_19.INIT0 = 16'hf555;
    defparam sub_2002_add_2_19.INIT1 = 16'hf555;
    defparam sub_2002_add_2_19.INJECT1_0 = "NO";
    defparam sub_2002_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27122), .COUT(n27123));
    defparam sub_2002_add_2_17.INIT0 = 16'hf555;
    defparam sub_2002_add_2_17.INIT1 = 16'hf555;
    defparam sub_2002_add_2_17.INJECT1_0 = "NO";
    defparam sub_2002_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27121), .COUT(n27122));
    defparam sub_2002_add_2_15.INIT0 = 16'hf555;
    defparam sub_2002_add_2_15.INIT1 = 16'hf555;
    defparam sub_2002_add_2_15.INJECT1_0 = "NO";
    defparam sub_2002_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27120), .COUT(n27121));
    defparam sub_2002_add_2_13.INIT0 = 16'hf555;
    defparam sub_2002_add_2_13.INIT1 = 16'hf555;
    defparam sub_2002_add_2_13.INJECT1_0 = "NO";
    defparam sub_2002_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27119), .COUT(n27120));
    defparam sub_2002_add_2_11.INIT0 = 16'hf555;
    defparam sub_2002_add_2_11.INIT1 = 16'hf555;
    defparam sub_2002_add_2_11.INJECT1_0 = "NO";
    defparam sub_2002_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27118), .COUT(n27119));
    defparam sub_2002_add_2_9.INIT0 = 16'hf555;
    defparam sub_2002_add_2_9.INIT1 = 16'hf555;
    defparam sub_2002_add_2_9.INJECT1_0 = "NO";
    defparam sub_2002_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27117), .COUT(n27118));
    defparam sub_2002_add_2_7.INIT0 = 16'hf555;
    defparam sub_2002_add_2_7.INIT1 = 16'hf555;
    defparam sub_2002_add_2_7.INJECT1_0 = "NO";
    defparam sub_2002_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27116), .COUT(n27117));
    defparam sub_2002_add_2_5.INIT0 = 16'hf555;
    defparam sub_2002_add_2_5.INIT1 = 16'hf555;
    defparam sub_2002_add_2_5.INJECT1_0 = "NO";
    defparam sub_2002_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27115), .COUT(n27116));
    defparam sub_2002_add_2_3.INIT0 = 16'hf555;
    defparam sub_2002_add_2_3.INIT1 = 16'hf555;
    defparam sub_2002_add_2_3.INJECT1_0 = "NO";
    defparam sub_2002_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2002_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27115));
    defparam sub_2002_add_2_1.INIT0 = 16'h0000;
    defparam sub_2002_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2002_add_2_1.INJECT1_0 = "NO";
    defparam sub_2002_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27298), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27297), .COUT(n27298), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27296), .COUT(n27297), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27295), .COUT(n27296), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27294), .COUT(n27295), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27293), .COUT(n27294), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27292), .COUT(n27293), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27291), .COUT(n27292), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27290), .COUT(n27291), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27289), .COUT(n27290), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27288), .COUT(n27289), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27287), .COUT(n27288), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27402), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_33.INIT1 = 16'h0000;
    defparam count_2579_add_4_33.INJECT1_0 = "NO";
    defparam count_2579_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27286), .COUT(n27287), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27285), .COUT(n27286), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27401), .COUT(n27402), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_31.INJECT1_0 = "NO";
    defparam count_2579_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27284), .COUT(n27285), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27400), .COUT(n27401), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_29.INJECT1_0 = "NO";
    defparam count_2579_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27399), .COUT(n27400), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_27.INJECT1_0 = "NO";
    defparam count_2579_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27398), .COUT(n27399), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_25.INJECT1_0 = "NO";
    defparam count_2579_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27283), .COUT(n27284), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27283), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27397), .COUT(n27398), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_23.INJECT1_0 = "NO";
    defparam count_2579_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27396), .COUT(n27397), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_21.INJECT1_0 = "NO";
    defparam count_2579_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27395), .COUT(n27396), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_19.INJECT1_0 = "NO";
    defparam count_2579_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27394), .COUT(n27395), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_17.INJECT1_0 = "NO";
    defparam count_2579_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27393), .COUT(n27394), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_15.INJECT1_0 = "NO";
    defparam count_2579_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27392), .COUT(n27393), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_13.INJECT1_0 = "NO";
    defparam count_2579_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27391), .COUT(n27392), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_11.INJECT1_0 = "NO";
    defparam count_2579_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27390), .COUT(n27391), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_9.INJECT1_0 = "NO";
    defparam count_2579_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27389), .COUT(n27390), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_7.INJECT1_0 = "NO";
    defparam count_2579_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27388), .COUT(n27389), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_5.INJECT1_0 = "NO";
    defparam count_2579_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27387), .COUT(n27388), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2579_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2579_add_4_3.INJECT1_0 = "NO";
    defparam count_2579_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2579_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27387), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579_add_4_1.INIT0 = 16'hF000;
    defparam count_2579_add_4_1.INIT1 = 16'h0555;
    defparam count_2579_add_4_1.INJECT1_0 = "NO";
    defparam count_2579_add_4_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31693), .CD(n16110), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31693), .PD(n16110), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1S3IX count_2579__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i1.GSR = "ENABLED";
    FD1S3IX count_2579__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i2.GSR = "ENABLED";
    FD1S3IX count_2579__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i3.GSR = "ENABLED";
    FD1S3IX count_2579__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i4.GSR = "ENABLED";
    FD1S3IX count_2579__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i5.GSR = "ENABLED";
    FD1S3IX count_2579__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i6.GSR = "ENABLED";
    FD1S3IX count_2579__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i7.GSR = "ENABLED";
    FD1S3IX count_2579__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i8.GSR = "ENABLED";
    FD1S3IX count_2579__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i9.GSR = "ENABLED";
    FD1S3IX count_2579__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i10.GSR = "ENABLED";
    FD1S3IX count_2579__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i11.GSR = "ENABLED";
    FD1S3IX count_2579__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i12.GSR = "ENABLED";
    FD1S3IX count_2579__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i13.GSR = "ENABLED";
    FD1S3IX count_2579__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i14.GSR = "ENABLED";
    FD1S3IX count_2579__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i15.GSR = "ENABLED";
    FD1S3IX count_2579__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i16.GSR = "ENABLED";
    FD1S3IX count_2579__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i17.GSR = "ENABLED";
    FD1S3IX count_2579__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i18.GSR = "ENABLED";
    FD1S3IX count_2579__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i19.GSR = "ENABLED";
    FD1S3IX count_2579__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i20.GSR = "ENABLED";
    FD1S3IX count_2579__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i21.GSR = "ENABLED";
    FD1S3IX count_2579__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i22.GSR = "ENABLED";
    FD1S3IX count_2579__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i23.GSR = "ENABLED";
    FD1S3IX count_2579__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i24.GSR = "ENABLED";
    FD1S3IX count_2579__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i25.GSR = "ENABLED";
    FD1S3IX count_2579__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i26.GSR = "ENABLED";
    FD1S3IX count_2579__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i27.GSR = "ENABLED";
    FD1S3IX count_2579__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i28.GSR = "ENABLED";
    FD1S3IX count_2579__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i29.GSR = "ENABLED";
    FD1S3IX count_2579__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i30.GSR = "ENABLED";
    FD1S3IX count_2579__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31693), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2579__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module SabertoothSerialPeripheral
//

module SabertoothSerialPeripheral (debug_c_c, n13476, n31699, n33451, 
            \databus[6] , \databus[5] , \databus[4] , \databus[3] , 
            \databus[2] , \register[1][1] , \databus[1] , \databus[0] , 
            \register[0] , n22093, n31698, \register[0][1] , \read_size[0] , 
            n106, n33450, \select[2] , n31867, n33447, \register_addr[0] , 
            n31832, n21959, n31796, n21892, n31818, rw, n5, n5_adj_5, 
            n5_adj_6, n5_adj_7, n5_adj_8, n5_adj_9, n5_adj_10, n5_adj_11, 
            \state[0] , n17748, n17735, n17753, n17745, GND_net, 
            n31695, \state[1] , n27884, n31, n21729, n31797, n19, 
            n9848, n7450, n44, n88, n42, n86, n45, n89, n43, 
            n87, \state[2] , n8110, select_clk, \reset_count[14] , 
            \reset_count[12] , \reset_count[13] , n31783, n31751, n24311, 
            n29370, n31784, \state[3] , n24417, n33449, n33453, 
            n33455, n31237, \reset_count[0] , \reset_count[3] , \reset_count[2] , 
            \reset_count[1] , n29966, n7485, n241, n29, \reset_count[5] , 
            \reset_count[6] , \reset_count[4] , \reset_count[11] , \reset_count[8] , 
            \reset_count[7] , n14424, n33448, \databus[7] , n31779, 
            n191, n31715, n9093, prev_select, n31774, \select[4] , 
            n2669, n28845, n33452, n31739, \register_addr[1] , n610, 
            n608, \register_addr[4] , prev_select_adj_12, n31763, n13671, 
            prev_select_adj_13, n14194, n579, motor_pwm_l_c) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n13476;
    input n31699;
    output n33451;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    output \register[1][1] ;
    input \databus[1] ;
    input \databus[0] ;
    output [7:0]\register[0] ;
    input n22093;
    input n31698;
    output \register[0][1] ;
    output \read_size[0] ;
    input n106;
    output n33450;
    input \select[2] ;
    output n31867;
    output n33447;
    input \register_addr[0] ;
    input n31832;
    output n21959;
    input n31796;
    output n21892;
    output n31818;
    input rw;
    output n5;
    output n5_adj_5;
    output n5_adj_6;
    output n5_adj_7;
    output n5_adj_8;
    output n5_adj_9;
    output n5_adj_10;
    output n5_adj_11;
    output \state[0] ;
    input n17748;
    input n17735;
    input n17753;
    input n17745;
    input GND_net;
    input n31695;
    output \state[1] ;
    input n27884;
    output n31;
    input n21729;
    input n31797;
    input n19;
    output n9848;
    input n7450;
    output n44;
    output n88;
    output n42;
    output n86;
    output n45;
    output n89;
    output n43;
    output n87;
    output \state[2] ;
    output n8110;
    output select_clk;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input \reset_count[13] ;
    output n31783;
    output n31751;
    input n24311;
    input n29370;
    output n31784;
    output \state[3] ;
    output n24417;
    output n33449;
    output n33453;
    output n33455;
    output n31237;
    input \reset_count[0] ;
    input \reset_count[3] ;
    input \reset_count[2] ;
    input \reset_count[1] ;
    output n29966;
    input n7485;
    output n241;
    output n29;
    input \reset_count[5] ;
    input \reset_count[6] ;
    input \reset_count[4] ;
    input \reset_count[11] ;
    input \reset_count[8] ;
    input \reset_count[7] ;
    input n14424;
    output n33448;
    input \databus[7] ;
    input n31779;
    input n191;
    input n31715;
    output n9093;
    input prev_select;
    input n31774;
    input \select[4] ;
    output n2669;
    input n28845;
    output n33452;
    input n31739;
    input \register_addr[1] ;
    output n610;
    output n608;
    input \register_addr[4] ;
    input prev_select_adj_12;
    input n31763;
    output n13671;
    input prev_select_adj_13;
    output n14194;
    output n579;
    output motor_pwm_l_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [15:0]n281;
    wire [7:0]\register[0]_c ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n2631, prev_select_c;
    wire [7:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(92[12:22])
    
    wire n9079;
    wire [7:0]n28;
    wire [31:0]n59;
    
    wire n31721, n27829, n21862, n27735, n21741;
    wire [31:0]n15;
    
    wire n21850, n27739;
    wire [7:0]n5984;
    
    FD1P3AX register_0__i16 (.D(n281[15]), .SP(n13476), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n31699), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n31699), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n31699), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n31699), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n31699), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n31699), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[1][1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n31699), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n281[15]), .SP(n22093), .CK(debug_c_c), 
            .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n31698), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[0]_c [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n31698), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[0]_c [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n31698), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[0]_c [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n31698), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[0]_c [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n31698), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[0]_c [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n31698), .PD(n33451), 
            .CK(debug_c_c), .Q(\register[0][1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i2.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n106), .SP(n2631), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n31698), .PD(n33450), 
            .CK(debug_c_c), .Q(\register[0]_c [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam prev_select_138.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n28[0]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_444 (.A(\select[2] ), .B(prev_select_c), .Z(n31867)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_rep_444.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\select[2] ), .B(prev_select_c), .C(n33447), 
         .Z(n2631)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 mux_1861_Mux_3_i1_3_lut (.A(\register[0]_c [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n28[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1861_Mux_4_i1_3_lut (.A(\register[0]_c [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n28[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1861_Mux_5_i1_3_lut (.A(\register[0]_c [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n28[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1861_Mux_6_i1_3_lut (.A(\register[0]_c [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n28[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1861_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n28[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 i15312_4_lut_4_lut (.A(\register[1][1] ), .B(n31832), .C(n21959), 
         .D(\register[1] [2]), .Z(n59[1])) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i15312_4_lut_4_lut.init = 16'hf1e2;
    LUT4 i23221_3_lut_4_lut_4_lut (.A(\register[1] [7]), .B(n31832), .C(n31796), 
         .D(n31721), .Z(n27829)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i23221_3_lut_4_lut_4_lut.init = 16'hfdff;
    LUT4 i1_4_lut_4_lut (.A(\register[1] [7]), .B(n31832), .C(n21862), 
         .D(n27735), .Z(n21959)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i1_4_lut_4_lut.init = 16'h2000;
    LUT4 i23196_3_lut_3_lut_4_lut (.A(\register[0][1] ), .B(n31832), .C(n21892), 
         .D(n31818), .Z(n21741)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i23196_3_lut_3_lut_4_lut.init = 16'h00f1;
    LUT4 i15305_4_lut_4_lut (.A(\register[0][1] ), .B(n31832), .C(n21892), 
         .D(\register[0]_c [2]), .Z(n15[1])) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i15305_4_lut_4_lut.init = 16'hf1e2;
    LUT4 i1_4_lut_4_lut_adj_9 (.A(\register[0] [7]), .B(n31832), .C(n21850), 
         .D(n27739), .Z(n21892)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i1_4_lut_4_lut_adj_9.init = 16'h2000;
    FD1P3IX read_value__i3 (.D(n28[3]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n28[4]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n28[5]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n28[6]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n28[7]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 mux_1861_Mux_2_i1_3_lut (.A(\register[0]_c [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n5984[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1861_Mux_1_i1_3_lut (.A(\register[0][1] ), .B(\register[1][1] ), 
         .C(\register_addr[0] ), .Z(n5984[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 Select_4198_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[0]), 
         .Z(n5)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4198_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4197_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[1]), 
         .Z(n5_adj_5)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4197_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4196_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[2]), 
         .Z(n5_adj_6)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4196_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4195_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[3]), 
         .Z(n5_adj_7)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4195_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4194_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[4]), 
         .Z(n5_adj_8)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4194_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4193_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[5]), 
         .Z(n5_adj_9)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4193_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4192_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[6]), 
         .Z(n5_adj_10)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4192_i5_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_4191_i5_2_lut_3_lut (.A(\select[2] ), .B(rw), .C(read_value[7]), 
         .Z(n5_adj_11)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam Select_4191_i5_2_lut_3_lut.init = 16'h8080;
    FD1P3IX read_value__i2 (.D(n5984[2]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n5984[1]), .SP(n2631), .CD(n9079), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=508, LSE_RLINE=516 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1861_Mux_0_i1_3_lut (.A(\register[0]_c [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n28[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1861_Mux_0_i1_3_lut.init = 16'hcaca;
    SabertoothSerial sserial (.\state[0] (\state[0] ), .n17748(n17748), 
            .n17735(n17735), .n17753(n17753), .n17745(n17745), .debug_c_c(debug_c_c), 
            .GND_net(GND_net), .n31695(n31695), .\register[1] ({\register[1] [7:2], 
            \register[1][1] , \register[1] [0]}), .\register[0] ({\register[0] [7], 
            \register[0]_c [6:2], \register[0][1] , \register[0]_c [0]}), 
            .n46(n15[1]), .n90(n59[1]), .\state[1] (\state[1] ), .n21862(n21862), 
            .n31818(n31818), .n27829(n27829), .n27884(n27884), .n31(n31), 
            .n21729(n21729), .n21741(n21741), .n31796(n31796), .n31797(n31797), 
            .n19(n19), .n31832(n31832), .n9848(n9848), .n7450(n7450), 
            .n44(n44), .n88(n88), .n42(n42), .n86(n86), .n31721(n31721), 
            .n45(n45), .n89(n89), .n43(n43), .n27739(n27739), .n21850(n21850), 
            .n87(n87), .n27735(n27735), .n33450(n33450), .\state[2] (\state[2] ), 
            .n33447(n33447), .n8110(n8110), .select_clk(select_clk), .\reset_count[14] (\reset_count[14] ), 
            .\reset_count[12] (\reset_count[12] ), .\reset_count[13] (\reset_count[13] ), 
            .n31783(n31783), .n31751(n31751), .n24311(n24311), .n29370(n29370), 
            .n31784(n31784), .\state[3] (\state[3] ), .n24417(n24417), 
            .n33449(n33449), .n33453(n33453), .n33455(n33455), .n31237(n31237), 
            .n33451(n33451), .\reset_count[0] (\reset_count[0] ), .\reset_count[3] (\reset_count[3] ), 
            .\reset_count[2] (\reset_count[2] ), .\reset_count[1] (\reset_count[1] ), 
            .n29966(n29966), .n7485(n7485), .n241(n241), .n29(n29), 
            .\reset_count[5] (\reset_count[5] ), .\reset_count[6] (\reset_count[6] ), 
            .\reset_count[4] (\reset_count[4] ), .\reset_count[11] (\reset_count[11] ), 
            .\reset_count[8] (\reset_count[8] ), .\reset_count[7] (\reset_count[7] ), 
            .n14424(n14424), .n33448(n33448), .\databus[7] (\databus[7] ), 
            .n282(n281[15]), .n31779(n31779), .n191(n191), .n31715(n31715), 
            .n9093(n9093), .prev_select(prev_select), .n31774(n31774), 
            .\select[4] (\select[4] ), .n2669(n2669), .n28845(n28845), 
            .n33452(n33452), .n31867(n31867), .n31739(n31739), .\register_addr[1] (\register_addr[1] ), 
            .n9079(n9079), .\databus[2] (\databus[2] ), .n610(n610), .\databus[4] (\databus[4] ), 
            .n608(n608), .\register_addr[4] (\register_addr[4] ), .prev_select_adj_3(prev_select_adj_12), 
            .n31763(n31763), .n13671(n13671), .prev_select_adj_4(prev_select_adj_13), 
            .n14194(n14194), .\databus[0] (\databus[0] ), .n579(n579), 
            .motor_pwm_l_c(motor_pwm_l_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(142[19] 147[34])
    
endmodule
//
// Verilog Description of module SabertoothSerial
//

module SabertoothSerial (\state[0] , n17748, n17735, n17753, n17745, 
            debug_c_c, GND_net, n31695, \register[1] , \register[0] , 
            n46, n90, \state[1] , n21862, n31818, n27829, n27884, 
            n31, n21729, n21741, n31796, n31797, n19, n31832, 
            n9848, n7450, n44, n88, n42, n86, n31721, n45, n89, 
            n43, n27739, n21850, n87, n27735, n33450, \state[2] , 
            n33447, n8110, select_clk, \reset_count[14] , \reset_count[12] , 
            \reset_count[13] , n31783, n31751, n24311, n29370, n31784, 
            \state[3] , n24417, n33449, n33453, n33455, n31237, 
            n33451, \reset_count[0] , \reset_count[3] , \reset_count[2] , 
            \reset_count[1] , n29966, n7485, n241, n29, \reset_count[5] , 
            \reset_count[6] , \reset_count[4] , \reset_count[11] , \reset_count[8] , 
            \reset_count[7] , n14424, n33448, \databus[7] , n282, 
            n31779, n191, n31715, n9093, prev_select, n31774, \select[4] , 
            n2669, n28845, n33452, n31867, n31739, \register_addr[1] , 
            n9079, \databus[2] , n610, \databus[4] , n608, \register_addr[4] , 
            prev_select_adj_3, n31763, n13671, prev_select_adj_4, n14194, 
            \databus[0] , n579, motor_pwm_l_c) /* synthesis syn_module_defined=1 */ ;
    output \state[0] ;
    input n17748;
    input n17735;
    input n17753;
    input n17745;
    input debug_c_c;
    input GND_net;
    input n31695;
    input [7:0]\register[1] ;
    input [7:0]\register[0] ;
    input n46;
    input n90;
    output \state[1] ;
    output n21862;
    output n31818;
    input n27829;
    input n27884;
    output n31;
    input n21729;
    input n21741;
    input n31796;
    input n31797;
    input n19;
    input n31832;
    output n9848;
    input n7450;
    output n44;
    output n88;
    output n42;
    output n86;
    output n31721;
    output n45;
    output n89;
    output n43;
    output n27739;
    output n21850;
    output n87;
    output n27735;
    output n33450;
    output \state[2] ;
    output n33447;
    output n8110;
    output select_clk;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input \reset_count[13] ;
    output n31783;
    output n31751;
    input n24311;
    input n29370;
    output n31784;
    output \state[3] ;
    output n24417;
    output n33449;
    output n33453;
    output n33455;
    output n31237;
    output n33451;
    input \reset_count[0] ;
    input \reset_count[3] ;
    input \reset_count[2] ;
    input \reset_count[1] ;
    output n29966;
    input n7485;
    output n241;
    output n29;
    input \reset_count[5] ;
    input \reset_count[6] ;
    input \reset_count[4] ;
    input \reset_count[11] ;
    input \reset_count[8] ;
    input \reset_count[7] ;
    input n14424;
    output n33448;
    input \databus[7] ;
    output n282;
    input n31779;
    input n191;
    input n31715;
    output n9093;
    input prev_select;
    input n31774;
    input \select[4] ;
    output n2669;
    input n28845;
    output n33452;
    input n31867;
    input n31739;
    input \register_addr[1] ;
    output n9079;
    input \databus[2] ;
    output n610;
    input \databus[4] ;
    output n608;
    input \register_addr[4] ;
    input prev_select_adj_3;
    input n31763;
    output n13671;
    input prev_select_adj_4;
    output n14194;
    input \databus[0] ;
    output n579;
    output motor_pwm_l_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n31848;
    wire [7:0]n5293;
    wire [3:0]n16;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(16[12:19])
    
    wire n21835, n31819, n31742, n31820, n31743, n33439, n976, 
        n31696, n31775, n31799, n31800, n31776, n7, n29_c, n26, 
        n107;
    
    LUT4 i3840_1_lut_rep_425 (.A(\state[0] ), .Z(n31848)) /* synthesis lut_function=(!(A)) */ ;
    defparam i3840_1_lut_rep_425.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(\state[0] ), .B(n17748), .Z(n5293[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_4 (.A(\state[0] ), .B(n17735), .Z(n5293[3])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_4.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_5 (.A(\state[0] ), .B(n17753), .Z(n5293[4])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_5.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_6 (.A(\state[0] ), .B(n17745), .Z(n5293[5])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_6.init = 16'h4444;
    FD1S3IX state__i0 (.D(n16[0]), .CK(debug_c_c), .CD(GND_net), .Q(\state[0] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n21835), .SP(n31695), .CK(debug_c_c), .Q(tx_data[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    LUT4 i6000_2_lut_rep_319_3_lut_4_lut (.A(\register[1] [3]), .B(n31819), 
         .C(\register[1] [5]), .D(\register[1] [4]), .Z(n31742)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6000_2_lut_rep_319_3_lut_4_lut.init = 16'h8000;
    LUT4 i5940_2_lut_rep_320_3_lut_4_lut (.A(\register[0] [3]), .B(n31820), 
         .C(\register[0] [5]), .D(\register[0] [4]), .Z(n31743)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5940_2_lut_rep_320_3_lut_4_lut.init = 16'h8000;
    LUT4 n46_bdd_4_lut (.A(n46), .B(n90), .C(\state[1] ), .D(\state[0] ), 
         .Z(n33439)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n46_bdd_4_lut.init = 16'h00ca;
    FD1P3IX send_27 (.D(n31848), .SP(n31696), .CD(GND_net), .CK(debug_c_c), 
            .Q(n976));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam send_27.GSR = "ENABLED";
    LUT4 i14983_2_lut (.A(\register[1] [0]), .B(\register[1] [4]), .Z(n21862)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14983_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_395 (.A(\state[0] ), .B(\state[1] ), .Z(n31818)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_395.init = 16'heeee;
    LUT4 i5103_2_lut_rep_396 (.A(\register[1] [2]), .B(\register[1] [1]), 
         .Z(n31819)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5103_2_lut_rep_396.init = 16'h8888;
    LUT4 i5998_2_lut_rep_352_3_lut_4_lut (.A(\register[1] [2]), .B(\register[1] [1]), 
         .C(\register[1] [4]), .D(\register[1] [3]), .Z(n31775)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5998_2_lut_rep_352_3_lut_4_lut.init = 16'h8000;
    LUT4 i5108_2_lut_rep_376_3_lut (.A(\register[1] [2]), .B(\register[1] [1]), 
         .C(\register[1] [3]), .Z(n31799)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5108_2_lut_rep_376_3_lut.init = 16'h8080;
    LUT4 i4540_2_lut_rep_397 (.A(\register[0] [2]), .B(\register[0] [1]), 
         .Z(n31820)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4540_2_lut_rep_397.init = 16'h8888;
    LUT4 i4562_2_lut_rep_377_3_lut (.A(\register[0] [2]), .B(\register[0] [1]), 
         .C(\register[0] [3]), .Z(n31800)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i4562_2_lut_rep_377_3_lut.init = 16'h8080;
    LUT4 i5898_2_lut_rep_353_3_lut_4_lut (.A(\register[0] [2]), .B(\register[0] [1]), 
         .C(\register[0] [4]), .D(\register[0] [3]), .Z(n31776)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5898_2_lut_rep_353_3_lut_4_lut.init = 16'h8000;
    PFUMX mux_1794_i8 (.BLUT(n27829), .ALUT(n27884), .C0(n7), .Z(n5293[7]));
    PFUMX i44 (.BLUT(n29_c), .ALUT(n26), .C0(\state[1] ), .Z(n31));
    PFUMX mux_1794_i1 (.BLUT(n21729), .ALUT(n21741), .C0(n7), .Z(n21835));
    FD1P3AX tx_data_i0_i1 (.D(n33439), .SP(n31695), .CK(debug_c_c), .Q(tx_data[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(\register[1] [6]), .B(n31742), .C(\register[1] [7]), 
         .D(n31796), .Z(n26)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A (C+(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0087;
    LUT4 i1_3_lut_4_lut_adj_7 (.A(\register[0] [6]), .B(n31743), .C(\register[0] [7]), 
         .D(n31797), .Z(n29_c)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_7.init = 16'h0087;
    FD1P3AX tx_data_i0_i2 (.D(n5293[2]), .SP(n31695), .CK(debug_c_c), 
            .Q(tx_data[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n5293[3]), .SP(n31695), .CK(debug_c_c), 
            .Q(tx_data[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n5293[4]), .SP(n31695), .CK(debug_c_c), 
            .Q(tx_data[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i5 (.D(n5293[5]), .SP(n31695), .CK(debug_c_c), 
            .Q(tx_data[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i6 (.D(n19), .SP(n31695), .CK(debug_c_c), .Q(tx_data[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i7 (.D(n5293[7]), .SP(n31695), .CK(debug_c_c), 
            .Q(tx_data[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i15446_2_lut_3_lut_4_lut (.A(\register[0] [5]), .B(n31776), .C(n31832), 
         .D(\register[0] [6]), .Z(n9848)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i15446_2_lut_3_lut_4_lut.init = 16'hf8f0;
    FD1P3IX state__i1 (.D(n7450), .SP(n31696), .CD(GND_net), .CK(debug_c_c), 
            .Q(\state[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 i15307_4_lut (.A(\register[0] [4]), .B(n31797), .C(n31832), .D(n31800), 
         .Z(n44)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(37[20:57])
    defparam i15307_4_lut.init = 16'hcdce;
    LUT4 i15314_4_lut (.A(\register[1] [4]), .B(n31796), .C(n31832), .D(n31799), 
         .Z(n88)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i15314_4_lut.init = 16'hcdce;
    LUT4 i15309_4_lut (.A(\register[0] [6]), .B(n31797), .C(n31832), .D(n31743), 
         .Z(n42)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(37[20:57])
    defparam i15309_4_lut.init = 16'hcdce;
    LUT4 i15316_4_lut (.A(\register[1] [6]), .B(n31796), .C(n31832), .D(n31742), 
         .Z(n86)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i15316_4_lut.init = 16'hcdce;
    LUT4 i6014_2_lut_rep_298_3_lut_4_lut (.A(\register[1] [4]), .B(n31799), 
         .C(\register[1] [6]), .D(\register[1] [5]), .Z(n31721)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6014_2_lut_rep_298_3_lut_4_lut.init = 16'h8000;
    LUT4 i15306_4_lut (.A(\register[0] [3]), .B(n31797), .C(n31832), .D(n31820), 
         .Z(n45)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(37[20:57])
    defparam i15306_4_lut.init = 16'hcdce;
    LUT4 i15313_4_lut (.A(\register[1] [3]), .B(n31796), .C(n31832), .D(n31819), 
         .Z(n89)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i15313_4_lut.init = 16'hcdce;
    LUT4 i15308_4_lut (.A(\register[0] [5]), .B(n31797), .C(n31832), .D(n31776), 
         .Z(n43)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(37[20:57])
    defparam i15308_4_lut.init = 16'hcdce;
    LUT4 i1_2_lut (.A(\state[0] ), .B(\state[1] ), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i3_4_lut (.A(\register[0] [2]), .B(\register[0] [6]), .C(\register[0] [5]), 
         .D(\register[0] [3]), .Z(n27739)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i14969_2_lut (.A(\register[0] [0]), .B(\register[0] [4]), .Z(n21850)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14969_2_lut.init = 16'h8888;
    LUT4 i15315_4_lut (.A(\register[1] [5]), .B(n31796), .C(n31832), .D(n31775), 
         .Z(n87)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:59])
    defparam i15315_4_lut.init = 16'hcdce;
    LUT4 i3_4_lut_adj_8 (.A(\register[1] [2]), .B(\register[1] [6]), .C(\register[1] [5]), 
         .D(\register[1] [3]), .Z(n27735)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_8.init = 16'h8000;
    \UARTTransmitter(baud_div=1250)  sender (.n33450(n33450), .\state[2] (\state[2] ), 
            .n33447(n33447), .\state[0] (\state[0] ), .n8110(n8110), .select_clk(select_clk), 
            .n12(n16[0]), .\reset_count[14] (\reset_count[14] ), .\reset_count[12] (\reset_count[12] ), 
            .\reset_count[13] (\reset_count[13] ), .n31783(n31783), .n31751(n31751), 
            .n24311(n24311), .n29370(n29370), .n31784(n31784), .\state[3] (\state[3] ), 
            .n24417(n24417), .n976(n976), .n33449(n33449), .n33453(n33453), 
            .n33455(n33455), .n31237(n31237), .n33451(n33451), .tx_data({tx_data}), 
            .\reset_count[0] (\reset_count[0] ), .\reset_count[3] (\reset_count[3] ), 
            .\reset_count[2] (\reset_count[2] ), .\reset_count[1] (\reset_count[1] ), 
            .n29966(n29966), .n7485(n7485), .n241(n241), .n29(n29), 
            .\reset_count[5] (\reset_count[5] ), .\reset_count[6] (\reset_count[6] ), 
            .\reset_count[4] (\reset_count[4] ), .\reset_count[11] (\reset_count[11] ), 
            .\reset_count[8] (\reset_count[8] ), .\reset_count[7] (\reset_count[7] ), 
            .n14424(n14424), .n31696(n31696), .n33448(n33448), .n107(n107), 
            .\databus[7] (\databus[7] ), .n282(n282), .n31779(n31779), 
            .n191(n191), .n31715(n31715), .n9093(n9093), .prev_select(prev_select), 
            .n31774(n31774), .\select[4] (\select[4] ), .n2669(n2669), 
            .n28845(n28845), .n33452(n33452), .n31867(n31867), .n31739(n31739), 
            .\register_addr[1] (\register_addr[1] ), .n9079(n9079), .\databus[2] (\databus[2] ), 
            .n610(n610), .\databus[4] (\databus[4] ), .n608(n608), .\register_addr[4] (\register_addr[4] ), 
            .prev_select_adj_1(prev_select_adj_3), .n31763(n31763), .n13671(n13671), 
            .prev_select_adj_2(prev_select_adj_4), .n14194(n14194), .\databus[0] (\databus[0] ), 
            .n579(n579), .motor_pwm_l_c(motor_pwm_l_c), .GND_net(GND_net), 
            .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(63[26] 67[47])
    \ClockDividerP(factor=12000)  baud_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .select_clk(select_clk), .n107(n107), .n8110(n8110), .n33447(n33447)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(21[25] 23[48])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=1250) 
//

module \UARTTransmitter(baud_div=1250)  (n33450, \state[2] , n33447, \state[0] , 
            n8110, select_clk, n12, \reset_count[14] , \reset_count[12] , 
            \reset_count[13] , n31783, n31751, n24311, n29370, n31784, 
            \state[3] , n24417, n976, n33449, n33453, n33455, n31237, 
            n33451, tx_data, \reset_count[0] , \reset_count[3] , \reset_count[2] , 
            \reset_count[1] , n29966, n7485, n241, n29, \reset_count[5] , 
            \reset_count[6] , \reset_count[4] , \reset_count[11] , \reset_count[8] , 
            \reset_count[7] , n14424, n31696, n33448, n107, \databus[7] , 
            n282, n31779, n191, n31715, n9093, prev_select, n31774, 
            \select[4] , n2669, n28845, n33452, n31867, n31739, 
            \register_addr[1] , n9079, \databus[2] , n610, \databus[4] , 
            n608, \register_addr[4] , prev_select_adj_1, n31763, n13671, 
            prev_select_adj_2, n14194, \databus[0] , n579, motor_pwm_l_c, 
            GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    output n33450;
    output \state[2] ;
    output n33447;
    input \state[0] ;
    input n8110;
    input select_clk;
    output n12;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input \reset_count[13] ;
    output n31783;
    output n31751;
    input n24311;
    input n29370;
    output n31784;
    output \state[3] ;
    output n24417;
    input n976;
    output n33449;
    output n33453;
    output n33455;
    output n31237;
    output n33451;
    input [7:0]tx_data;
    input \reset_count[0] ;
    input \reset_count[3] ;
    input \reset_count[2] ;
    input \reset_count[1] ;
    output n29966;
    input n7485;
    output n241;
    output n29;
    input \reset_count[5] ;
    input \reset_count[6] ;
    input \reset_count[4] ;
    input \reset_count[11] ;
    input \reset_count[8] ;
    input \reset_count[7] ;
    input n14424;
    output n31696;
    output n33448;
    output n107;
    input \databus[7] ;
    output n282;
    input n31779;
    input n191;
    input n31715;
    output n9093;
    input prev_select;
    input n31774;
    input \select[4] ;
    output n2669;
    input n28845;
    output n33452;
    input n31867;
    input n31739;
    input \register_addr[1] ;
    output n9079;
    input \databus[2] ;
    output n610;
    input \databus[4] ;
    output n608;
    input \register_addr[4] ;
    input prev_select_adj_1;
    input n31763;
    output n13671;
    input prev_select_adj_2;
    output n14194;
    input \databus[0] ;
    output n579;
    output motor_pwm_l_c;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n30695, n2, n30043, n7;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n10, n27737, n238, n27753, n30041, n30042, n30694, n30693, 
        n29942, n8999, n27734, n21231, n29430, n104, n30832;
    
    FD1S3IX state__i0 (.D(n30695), .CK(bclk), .CD(n33450), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n30043), .C(\state[2] ), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15347_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15347_4_lut.init = 16'hfcee;
    LUT4 i1_3_lut_4_lut_4_lut_3_lut_4_lut (.A(n33447), .B(\state[0] ), .C(n8110), 
         .D(select_clk), .Z(n12)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hcc9c;
    LUT4 i1_4_lut_rep_360 (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n27737), .Z(n31783)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i1_4_lut_rep_360.init = 16'hfaea;
    LUT4 i55_1_lut_rep_328_4_lut (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n27737), .Z(n31751)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i55_1_lut_rep_328_4_lut.init = 16'h0515;
    LUT4 i23252_4_lut_rep_361 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n31784)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_361.init = 16'h575f;
    LUT4 i2_4_lut (.A(\state[2] ), .B(n33447), .C(\state[3] ), .D(n24417), 
         .Z(n27753)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    defparam i2_4_lut.init = 16'h1210;
    LUT4 i1_2_lut (.A(state[1]), .B(state[0]), .Z(n24417)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i23252_4_lut_rep_452 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n33447)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_452.init = 16'h575f;
    LUT4 i22888_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n30041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22888_3_lut.init = 16'hcaca;
    LUT4 i22889_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n30042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22889_3_lut.init = 16'hcaca;
    LUT4 n976_bdd_4_lut_23522 (.A(n976), .B(state[1]), .C(\state[3] ), 
         .D(state[0]), .Z(n30694)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam n976_bdd_4_lut_23522.init = 16'h80fe;
    LUT4 i23252_4_lut_rep_454 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n33449)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_454.init = 16'h575f;
    LUT4 n976_bdd_2_lut_23521 (.A(\state[3] ), .B(state[0]), .Z(n30693)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam n976_bdd_2_lut_23521.init = 16'h1111;
    LUT4 i23252_4_lut_rep_458 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n33453)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_458.init = 16'h575f;
    LUT4 i55_1_lut_rep_460 (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n27737), .Z(n33455)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i55_1_lut_rep_460.init = 16'h0515;
    LUT4 i23252_4_lut_rep_455 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n33450)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_455.init = 16'h575f;
    LUT4 i22792_2_lut_3_lut (.A(\state[2] ), .B(state[0]), .C(\state[3] ), 
         .Z(n29942)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22792_2_lut_3_lut.init = 16'hfefe;
    LUT4 n976_bdd_4_lut (.A(n976), .B(\state[3] ), .C(state[0]), .D(state[1]), 
         .Z(n31237)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam n976_bdd_4_lut.init = 16'h7ffe;
    LUT4 i23252_4_lut_rep_456 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n33451)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_456.init = 16'h575f;
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n8999), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 i22814_4_lut (.A(\reset_count[0] ), .B(\reset_count[3] ), .C(\reset_count[2] ), 
         .D(\reset_count[1] ), .Z(n29966)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22814_4_lut.init = 16'hfffe;
    LUT4 i14755_2_lut_2_lut (.A(n33447), .B(n7485), .Z(n241)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14755_2_lut_2_lut.init = 16'h4444;
    LUT4 i202_4_lut (.A(n29), .B(\reset_count[5] ), .C(\reset_count[6] ), 
         .D(\reset_count[4] ), .Z(n238)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i202_4_lut.init = 16'hfaea;
    LUT4 i2_4_lut_adj_1 (.A(n24311), .B(n27734), .C(\reset_count[11] ), 
         .D(\reset_count[8] ), .Z(n27737)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i2_4_lut_adj_1.init = 16'ha080;
    LUT4 i2_3_lut (.A(\reset_count[6] ), .B(\reset_count[7] ), .C(\reset_count[5] ), 
         .Z(n27734)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i1_4_lut (.A(n33447), .B(state[1]), .C(n21231), .D(state[0]), 
         .Z(n29430)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0104;
    LUT4 i14861_2_lut (.A(\state[2] ), .B(\state[3] ), .Z(n21231)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14861_2_lut.init = 16'h8888;
    LUT4 i20545_2_lut (.A(\reset_count[7] ), .B(\reset_count[8] ), .Z(n29)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    defparam i20545_2_lut.init = 16'heeee;
    FD1P3AX state__i3 (.D(n27753), .SP(n14424), .CK(bclk), .Q(\state[3] )) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_273_3_lut_3_lut (.A(n33447), .B(select_clk), .C(n8110), 
         .Z(n31696)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_273_3_lut_3_lut.init = 16'h1010;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(\state[3] ), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;
    LUT4 i23252_4_lut_rep_453 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n33448)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_453.init = 16'h575f;
    PFUMX i23349 (.BLUT(n30694), .ALUT(n30693), .C0(\state[2] ), .Z(n30695));
    PFUMX i22890 (.BLUT(n30041), .ALUT(n30042), .C0(state[1]), .Z(n30043));
    LUT4 i1_2_lut_2_lut (.A(n33447), .B(n8110), .Z(n107)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 state_3__bdd_4_lut (.A(\state[3] ), .B(\state[2] ), .C(state[0]), 
         .D(state[1]), .Z(n30832)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B+(C+(D))))) */ ;
    defparam state_3__bdd_4_lut.init = 16'h5776;
    LUT4 i15422_2_lut_2_lut (.A(n33447), .B(\databus[7] ), .Z(n282)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15422_2_lut_2_lut.init = 16'h4444;
    LUT4 i2_4_lut_4_lut (.A(n33447), .B(n31779), .C(n191), .D(n31715), 
         .Z(n9093)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C+!(D))))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h4500;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n33447), .B(prev_select), .C(n31774), 
         .D(\select[4] ), .Z(n2669)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    FD1P3AX state__i2 (.D(n28845), .SP(n14424), .CK(bclk), .Q(\state[2] )) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n29430), .SP(n14424), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 i23252_4_lut_rep_457 (.A(\reset_count[14] ), .B(n24311), .C(n29370), 
         .D(n238), .Z(n33452)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23252_4_lut_rep_457.init = 16'h575f;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n33447), .B(n31867), .C(n31739), .D(\register_addr[1] ), 
         .Z(n9079)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut.init = 16'h4440;
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n8999), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    LUT4 i15433_2_lut_2_lut (.A(n33447), .B(\databus[2] ), .Z(n610)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15433_2_lut_2_lut.init = 16'h4444;
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n8999), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n8999), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n8999), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n8999), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n8999), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n8999), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i15440_2_lut_2_lut (.A(n33447), .B(\databus[4] ), .Z(n608)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15440_2_lut_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_4_lut_4_lut_adj_2 (.A(n33447), .B(\register_addr[4] ), 
         .C(prev_select_adj_1), .D(n31763), .Z(n13671)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut_adj_2.init = 16'h0100;
    LUT4 i2_3_lut_4_lut_4_lut_adj_3 (.A(n33447), .B(prev_select_adj_2), 
         .C(\register_addr[4] ), .D(n31763), .Z(n14194)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut_adj_3.init = 16'h1000;
    LUT4 i4_4_lut (.A(n29942), .B(state[1]), .C(n976), .D(n33447), .Z(n8999)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i4_4_lut.init = 16'h0010;
    LUT4 i15028_2_lut_2_lut (.A(n33447), .B(\databus[0] ), .Z(n579)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15028_2_lut_2_lut.init = 16'h4444;
    FD1P3JX tx_35 (.D(n104), .SP(n30832), .PD(n33453), .CK(bclk), .Q(motor_pwm_l_c)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    \ClockDividerP(factor=1250)  baud_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .bclk(bclk)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=1250) 
//

module \ClockDividerP(factor=1250)  (GND_net, debug_c_c, bclk) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    output bclk;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    
    wire n27593;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n102;
    
    wire n27594, n27592, n27591, n27590, n27589, n27588, n27587, 
        n16108, n28243, n8, n39, n52, n48, n40, n31, n50, 
        n44, n32, n42, n46, n36, n8145, n27497, n27496, n27495, 
        n27494, n27493, n27492, n27491, n27490, n27489, n27488, 
        n27487, n27486, n27485, n27484, n27483, n27602, n27601, 
        n27600, n27599, n27598, n27597, n27596, n27595;
    
    CCU2D count_2585_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27593), .COUT(n27594), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_15.INJECT1_0 = "NO";
    defparam count_2585_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27592), .COUT(n27593), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_13.INJECT1_0 = "NO";
    defparam count_2585_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27591), .COUT(n27592), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_11.INJECT1_0 = "NO";
    defparam count_2585_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27590), .COUT(n27591), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_9.INJECT1_0 = "NO";
    defparam count_2585_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27589), .COUT(n27590), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_7.INJECT1_0 = "NO";
    defparam count_2585_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27588), .COUT(n27589), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_5.INJECT1_0 = "NO";
    defparam count_2585_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27587), .COUT(n27588), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_3.INJECT1_0 = "NO";
    defparam count_2585_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27587), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_1.INIT0 = 16'hF000;
    defparam count_2585_add_4_1.INIT1 = 16'h0555;
    defparam count_2585_add_4_1.INJECT1_0 = "NO";
    defparam count_2585_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2585__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i0.GSR = "ENABLED";
    LUT4 i23166_4_lut (.A(n28243), .B(count[5]), .C(n8), .D(count[0]), 
         .Z(n16108)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23166_4_lut.init = 16'h4000;
    LUT4 i26_4_lut (.A(n39), .B(n52), .C(n48), .D(n40), .Z(n28243)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i3_3_lut (.A(count[10]), .B(count[6]), .C(count[7]), .Z(n8)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3_3_lut.init = 16'h8080;
    LUT4 i12_2_lut (.A(count[30]), .B(count[13]), .Z(n39)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i12_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(n31), .B(n50), .C(n44), .D(n32), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(count[27]), .B(n42), .C(count[23]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(count[22]), .B(count[18]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i4_2_lut (.A(count[28]), .B(count[9]), .Z(n31)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(count[19]), .B(n46), .C(n36), .D(count[25]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(count[4]), .B(count[11]), .C(count[8]), .D(count[14]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[12]), .B(count[1]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[20]), .B(count[2]), .C(count[24]), .D(count[29]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(count[26]), .B(count[3]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i15_4_lut (.A(count[16]), .B(count[15]), .C(count[31]), .D(count[21]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_4_lut.init = 16'hfffe;
    FD1S3AX clk_o_14 (.D(n8145), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D add_20539_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27497), 
          .S1(n8145));
    defparam add_20539_32.INIT0 = 16'h5555;
    defparam add_20539_32.INIT1 = 16'h0000;
    defparam add_20539_32.INJECT1_0 = "NO";
    defparam add_20539_32.INJECT1_1 = "NO";
    CCU2D add_20539_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27496), .COUT(n27497));
    defparam add_20539_30.INIT0 = 16'h5555;
    defparam add_20539_30.INIT1 = 16'h5555;
    defparam add_20539_30.INJECT1_0 = "NO";
    defparam add_20539_30.INJECT1_1 = "NO";
    CCU2D add_20539_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27495), .COUT(n27496));
    defparam add_20539_28.INIT0 = 16'h5555;
    defparam add_20539_28.INIT1 = 16'h5555;
    defparam add_20539_28.INJECT1_0 = "NO";
    defparam add_20539_28.INJECT1_1 = "NO";
    CCU2D add_20539_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27494), .COUT(n27495));
    defparam add_20539_26.INIT0 = 16'h5555;
    defparam add_20539_26.INIT1 = 16'h5555;
    defparam add_20539_26.INJECT1_0 = "NO";
    defparam add_20539_26.INJECT1_1 = "NO";
    CCU2D add_20539_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27493), .COUT(n27494));
    defparam add_20539_24.INIT0 = 16'h5555;
    defparam add_20539_24.INIT1 = 16'h5555;
    defparam add_20539_24.INJECT1_0 = "NO";
    defparam add_20539_24.INJECT1_1 = "NO";
    CCU2D add_20539_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27492), .COUT(n27493));
    defparam add_20539_22.INIT0 = 16'h5555;
    defparam add_20539_22.INIT1 = 16'h5555;
    defparam add_20539_22.INJECT1_0 = "NO";
    defparam add_20539_22.INJECT1_1 = "NO";
    CCU2D add_20539_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27491), .COUT(n27492));
    defparam add_20539_20.INIT0 = 16'h5555;
    defparam add_20539_20.INIT1 = 16'h5555;
    defparam add_20539_20.INJECT1_0 = "NO";
    defparam add_20539_20.INJECT1_1 = "NO";
    CCU2D add_20539_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27490), .COUT(n27491));
    defparam add_20539_18.INIT0 = 16'h5555;
    defparam add_20539_18.INIT1 = 16'h5555;
    defparam add_20539_18.INJECT1_0 = "NO";
    defparam add_20539_18.INJECT1_1 = "NO";
    FD1S3IX count_2585__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i1.GSR = "ENABLED";
    CCU2D add_20539_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27489), .COUT(n27490));
    defparam add_20539_16.INIT0 = 16'h5555;
    defparam add_20539_16.INIT1 = 16'h5555;
    defparam add_20539_16.INJECT1_0 = "NO";
    defparam add_20539_16.INJECT1_1 = "NO";
    FD1S3IX count_2585__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i2.GSR = "ENABLED";
    FD1S3IX count_2585__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i3.GSR = "ENABLED";
    FD1S3IX count_2585__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i4.GSR = "ENABLED";
    FD1S3IX count_2585__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i5.GSR = "ENABLED";
    FD1S3IX count_2585__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i6.GSR = "ENABLED";
    FD1S3IX count_2585__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i7.GSR = "ENABLED";
    FD1S3IX count_2585__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i8.GSR = "ENABLED";
    FD1S3IX count_2585__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i9.GSR = "ENABLED";
    FD1S3IX count_2585__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i10.GSR = "ENABLED";
    FD1S3IX count_2585__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i11.GSR = "ENABLED";
    FD1S3IX count_2585__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i12.GSR = "ENABLED";
    FD1S3IX count_2585__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i13.GSR = "ENABLED";
    FD1S3IX count_2585__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i14.GSR = "ENABLED";
    FD1S3IX count_2585__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i15.GSR = "ENABLED";
    FD1S3IX count_2585__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i16.GSR = "ENABLED";
    FD1S3IX count_2585__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i17.GSR = "ENABLED";
    FD1S3IX count_2585__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i18.GSR = "ENABLED";
    FD1S3IX count_2585__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i19.GSR = "ENABLED";
    FD1S3IX count_2585__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i20.GSR = "ENABLED";
    FD1S3IX count_2585__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i21.GSR = "ENABLED";
    FD1S3IX count_2585__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i22.GSR = "ENABLED";
    FD1S3IX count_2585__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i23.GSR = "ENABLED";
    FD1S3IX count_2585__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i24.GSR = "ENABLED";
    FD1S3IX count_2585__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i25.GSR = "ENABLED";
    FD1S3IX count_2585__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i26.GSR = "ENABLED";
    FD1S3IX count_2585__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i27.GSR = "ENABLED";
    FD1S3IX count_2585__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i28.GSR = "ENABLED";
    FD1S3IX count_2585__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i29.GSR = "ENABLED";
    FD1S3IX count_2585__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i30.GSR = "ENABLED";
    FD1S3IX count_2585__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16108), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585__i31.GSR = "ENABLED";
    CCU2D add_20539_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27488), .COUT(n27489));
    defparam add_20539_14.INIT0 = 16'h5555;
    defparam add_20539_14.INIT1 = 16'h5555;
    defparam add_20539_14.INJECT1_0 = "NO";
    defparam add_20539_14.INJECT1_1 = "NO";
    CCU2D add_20539_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27487), .COUT(n27488));
    defparam add_20539_12.INIT0 = 16'h5555;
    defparam add_20539_12.INIT1 = 16'h5555;
    defparam add_20539_12.INJECT1_0 = "NO";
    defparam add_20539_12.INJECT1_1 = "NO";
    CCU2D add_20539_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27486), .COUT(n27487));
    defparam add_20539_10.INIT0 = 16'h5aaa;
    defparam add_20539_10.INIT1 = 16'h5555;
    defparam add_20539_10.INJECT1_0 = "NO";
    defparam add_20539_10.INJECT1_1 = "NO";
    CCU2D add_20539_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27485), 
          .COUT(n27486));
    defparam add_20539_8.INIT0 = 16'h5555;
    defparam add_20539_8.INIT1 = 16'h5555;
    defparam add_20539_8.INJECT1_0 = "NO";
    defparam add_20539_8.INJECT1_1 = "NO";
    CCU2D add_20539_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27484), 
          .COUT(n27485));
    defparam add_20539_6.INIT0 = 16'h5aaa;
    defparam add_20539_6.INIT1 = 16'h5aaa;
    defparam add_20539_6.INJECT1_0 = "NO";
    defparam add_20539_6.INJECT1_1 = "NO";
    CCU2D add_20539_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27483), 
          .COUT(n27484));
    defparam add_20539_4.INIT0 = 16'h5555;
    defparam add_20539_4.INIT1 = 16'h5aaa;
    defparam add_20539_4.INJECT1_0 = "NO";
    defparam add_20539_4.INJECT1_1 = "NO";
    CCU2D add_20539_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27483));
    defparam add_20539_2.INIT0 = 16'h1000;
    defparam add_20539_2.INIT1 = 16'h5555;
    defparam add_20539_2.INJECT1_0 = "NO";
    defparam add_20539_2.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27602), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_33.INIT1 = 16'h0000;
    defparam count_2585_add_4_33.INJECT1_0 = "NO";
    defparam count_2585_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27601), .COUT(n27602), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_31.INJECT1_0 = "NO";
    defparam count_2585_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27600), .COUT(n27601), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_29.INJECT1_0 = "NO";
    defparam count_2585_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27599), .COUT(n27600), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_27.INJECT1_0 = "NO";
    defparam count_2585_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27598), .COUT(n27599), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_25.INJECT1_0 = "NO";
    defparam count_2585_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27597), .COUT(n27598), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_23.INJECT1_0 = "NO";
    defparam count_2585_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27596), .COUT(n27597), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_21.INJECT1_0 = "NO";
    defparam count_2585_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27595), .COUT(n27596), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_19.INJECT1_0 = "NO";
    defparam count_2585_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2585_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27594), .COUT(n27595), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2585_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2585_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2585_add_4_17.INJECT1_0 = "NO";
    defparam count_2585_add_4_17.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000) 
//

module \ClockDividerP(factor=12000)  (GND_net, debug_c_c, select_clk, 
            n107, n8110, n33447) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    output select_clk;
    input n107;
    output n8110;
    input n33447;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27586;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n27585, n27584, n27583, n27582, n27581, n27580, n27579, 
        n27578, n27577, n27576, n27575, n27574, n27573, n27572, 
        n27571, n2770, n27510, n27509, n27508, n27507, n27506, 
        n27505, n27504, n27503, n27502, n27501, n27500, n27499, 
        n27498, n30137, n28239, n15, n20, n16, n27, n40, n36, 
        n28, n18, n38, n32, n34, n24;
    
    CCU2D count_2584_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27586), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_33.INIT1 = 16'h0000;
    defparam count_2584_add_4_33.INJECT1_0 = "NO";
    defparam count_2584_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27585), .COUT(n27586), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_31.INJECT1_0 = "NO";
    defparam count_2584_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27584), .COUT(n27585), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_29.INJECT1_0 = "NO";
    defparam count_2584_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27583), .COUT(n27584), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_27.INJECT1_0 = "NO";
    defparam count_2584_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27582), .COUT(n27583), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_25.INJECT1_0 = "NO";
    defparam count_2584_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27581), .COUT(n27582), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_23.INJECT1_0 = "NO";
    defparam count_2584_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27580), .COUT(n27581), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_21.INJECT1_0 = "NO";
    defparam count_2584_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27579), .COUT(n27580), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_19.INJECT1_0 = "NO";
    defparam count_2584_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27578), .COUT(n27579), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_17.INJECT1_0 = "NO";
    defparam count_2584_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27577), .COUT(n27578), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_15.INJECT1_0 = "NO";
    defparam count_2584_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27576), .COUT(n27577), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_13.INJECT1_0 = "NO";
    defparam count_2584_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27575), .COUT(n27576), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_11.INJECT1_0 = "NO";
    defparam count_2584_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27574), .COUT(n27575), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_9.INJECT1_0 = "NO";
    defparam count_2584_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27573), .COUT(n27574), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_7.INJECT1_0 = "NO";
    defparam count_2584_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27572), .COUT(n27573), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_5.INJECT1_0 = "NO";
    defparam count_2584_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27571), .COUT(n27572), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2584_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2584_add_4_3.INJECT1_0 = "NO";
    defparam count_2584_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2584_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27571), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584_add_4_1.INIT0 = 16'hF000;
    defparam count_2584_add_4_1.INIT1 = 16'h0555;
    defparam count_2584_add_4_1.INJECT1_0 = "NO";
    defparam count_2584_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2584__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2770), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i0.GSR = "ENABLED";
    FD1S3AX clk_o_14 (.D(n107), .CK(debug_c_c), .Q(select_clk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=25, LSE_RCOL=48, LSE_LLINE=21, LSE_RLINE=23 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D add_20538_28 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27510), 
          .S1(n8110));
    defparam add_20538_28.INIT0 = 16'h5555;
    defparam add_20538_28.INIT1 = 16'h0000;
    defparam add_20538_28.INJECT1_0 = "NO";
    defparam add_20538_28.INJECT1_1 = "NO";
    CCU2D add_20538_26 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27509), .COUT(n27510));
    defparam add_20538_26.INIT0 = 16'h5555;
    defparam add_20538_26.INIT1 = 16'h5555;
    defparam add_20538_26.INJECT1_0 = "NO";
    defparam add_20538_26.INJECT1_1 = "NO";
    CCU2D add_20538_24 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27508), .COUT(n27509));
    defparam add_20538_24.INIT0 = 16'h5555;
    defparam add_20538_24.INIT1 = 16'h5555;
    defparam add_20538_24.INJECT1_0 = "NO";
    defparam add_20538_24.INJECT1_1 = "NO";
    CCU2D add_20538_22 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27507), .COUT(n27508));
    defparam add_20538_22.INIT0 = 16'h5555;
    defparam add_20538_22.INIT1 = 16'h5555;
    defparam add_20538_22.INJECT1_0 = "NO";
    defparam add_20538_22.INJECT1_1 = "NO";
    CCU2D add_20538_20 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27506), .COUT(n27507));
    defparam add_20538_20.INIT0 = 16'h5555;
    defparam add_20538_20.INIT1 = 16'h5555;
    defparam add_20538_20.INJECT1_0 = "NO";
    defparam add_20538_20.INJECT1_1 = "NO";
    CCU2D add_20538_18 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27505), .COUT(n27506));
    defparam add_20538_18.INIT0 = 16'h5555;
    defparam add_20538_18.INIT1 = 16'h5555;
    defparam add_20538_18.INJECT1_0 = "NO";
    defparam add_20538_18.INJECT1_1 = "NO";
    CCU2D add_20538_16 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27504), .COUT(n27505));
    defparam add_20538_16.INIT0 = 16'h5555;
    defparam add_20538_16.INIT1 = 16'h5555;
    defparam add_20538_16.INJECT1_0 = "NO";
    defparam add_20538_16.INJECT1_1 = "NO";
    CCU2D add_20538_14 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27503), .COUT(n27504));
    defparam add_20538_14.INIT0 = 16'h5555;
    defparam add_20538_14.INIT1 = 16'h5555;
    defparam add_20538_14.INJECT1_0 = "NO";
    defparam add_20538_14.INJECT1_1 = "NO";
    CCU2D add_20538_12 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27502), .COUT(n27503));
    defparam add_20538_12.INIT0 = 16'h5555;
    defparam add_20538_12.INIT1 = 16'h5555;
    defparam add_20538_12.INJECT1_0 = "NO";
    defparam add_20538_12.INJECT1_1 = "NO";
    CCU2D add_20538_10 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27501), .COUT(n27502));
    defparam add_20538_10.INIT0 = 16'h5555;
    defparam add_20538_10.INIT1 = 16'h5555;
    defparam add_20538_10.INJECT1_0 = "NO";
    defparam add_20538_10.INJECT1_1 = "NO";
    CCU2D add_20538_8 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27500), .COUT(n27501));
    defparam add_20538_8.INIT0 = 16'h5555;
    defparam add_20538_8.INIT1 = 16'h5aaa;
    defparam add_20538_8.INJECT1_0 = "NO";
    defparam add_20538_8.INJECT1_1 = "NO";
    CCU2D add_20538_6 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27499), .COUT(n27500));
    defparam add_20538_6.INIT0 = 16'h5aaa;
    defparam add_20538_6.INIT1 = 16'h5aaa;
    defparam add_20538_6.INJECT1_0 = "NO";
    defparam add_20538_6.INJECT1_1 = "NO";
    CCU2D add_20538_4 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27498), 
          .COUT(n27499));
    defparam add_20538_4.INIT0 = 16'h5555;
    defparam add_20538_4.INIT1 = 16'h5aaa;
    defparam add_20538_4.INJECT1_0 = "NO";
    defparam add_20538_4.INJECT1_1 = "NO";
    CCU2D add_20538_2 (.A0(count[5]), .B0(count[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27498));
    defparam add_20538_2.INIT0 = 16'h7000;
    defparam add_20538_2.INIT1 = 16'h5aaa;
    defparam add_20538_2.INJECT1_0 = "NO";
    defparam add_20538_2.INJECT1_1 = "NO";
    LUT4 i23084_2_lut (.A(n30137), .B(n33447), .Z(n2770)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23084_2_lut.init = 16'heeee;
    LUT4 i23082_4_lut (.A(n28239), .B(n15), .C(n20), .D(n16), .Z(n30137)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i23082_4_lut.init = 16'h4000;
    LUT4 i20_4_lut (.A(n27), .B(n40), .C(n36), .D(n28), .Z(n28239)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[11]), .B(count[10]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(count[9]), .B(n18), .C(count[6]), .D(count[7]), 
         .Z(n20)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(count[1]), .B(count[4]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i6_2_lut (.A(count[28]), .B(count[12]), .Z(n27)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[5]), .B(n38), .C(n32), .D(count[20]), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(count[8]), .B(count[25]), .C(count[15]), .D(count[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[17]), .B(count[24]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i7_4_lut (.A(count[13]), .B(count[2]), .C(count[3]), .D(count[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i17_4_lut (.A(count[29]), .B(n34), .C(n24), .D(count[14]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(count[22]), .B(count[21]), .C(count[31]), .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(count[16]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[19]), .B(count[18]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    FD1S3IX count_2584__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2770), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i1.GSR = "ENABLED";
    FD1S3IX count_2584__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2770), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i2.GSR = "ENABLED";
    FD1S3IX count_2584__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2770), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i3.GSR = "ENABLED";
    FD1S3IX count_2584__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2770), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i4.GSR = "ENABLED";
    FD1S3IX count_2584__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2770), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i5.GSR = "ENABLED";
    FD1S3IX count_2584__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2770), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i6.GSR = "ENABLED";
    FD1S3IX count_2584__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2770), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i7.GSR = "ENABLED";
    FD1S3IX count_2584__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2770), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i8.GSR = "ENABLED";
    FD1S3IX count_2584__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2770), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i9.GSR = "ENABLED";
    FD1S3IX count_2584__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i10.GSR = "ENABLED";
    FD1S3IX count_2584__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i11.GSR = "ENABLED";
    FD1S3IX count_2584__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i12.GSR = "ENABLED";
    FD1S3IX count_2584__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i13.GSR = "ENABLED";
    FD1S3IX count_2584__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i14.GSR = "ENABLED";
    FD1S3IX count_2584__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i15.GSR = "ENABLED";
    FD1S3IX count_2584__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i16.GSR = "ENABLED";
    FD1S3IX count_2584__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i17.GSR = "ENABLED";
    FD1S3IX count_2584__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i18.GSR = "ENABLED";
    FD1S3IX count_2584__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i19.GSR = "ENABLED";
    FD1S3IX count_2584__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i20.GSR = "ENABLED";
    FD1S3IX count_2584__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i21.GSR = "ENABLED";
    FD1S3IX count_2584__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i22.GSR = "ENABLED";
    FD1S3IX count_2584__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i23.GSR = "ENABLED";
    FD1S3IX count_2584__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i24.GSR = "ENABLED";
    FD1S3IX count_2584__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i25.GSR = "ENABLED";
    FD1S3IX count_2584__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i26.GSR = "ENABLED";
    FD1S3IX count_2584__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i27.GSR = "ENABLED";
    FD1S3IX count_2584__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i28.GSR = "ENABLED";
    FD1S3IX count_2584__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i29.GSR = "ENABLED";
    FD1S3IX count_2584__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i30.GSR = "ENABLED";
    FD1S3IX count_2584__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2770), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2584__i31.GSR = "ENABLED";
    
endmodule
